`define PX 509'h136cf14c6c616b9ea31bd7eb68b8f08d1ca3e0019398e2d1e73054d0f3fa711f09da5ccd3ade6e68dc4ce3f375d535083f9434ac4a3b2f4bee6578e1bf6b3a33

`define PX_ 509'h1e865b392d85efd59d21ac99107fc69aee6e847c97f9bba4bb9ac32ec161f9c589428f2413a3287f37e786cfbe59ecaaecf885b245263b4b2d798abf9549878

`define PX3 509'hf9c25e546b0ada3ef77a25846a8f7b9bed60f720099ab5d4fbcfc6b1bce31e658b20ae8b86a0958f54ff3197e09f772e1f523f6019667e288b64789ccc20943

`define PY 509'hdcbf8519c6ed502ce81461020b9dd0e7e21ba5a0bbe0f864b03f6def88d71b967e5432476fc772c7a096d7218ee2541fb55bd9d37007684f07cfe55919d181a

`define PY_ 509'h7895eae62caf5992e6caca4d9070fe84d690def515a6f05e7e60a24e7831f01fa89429b051c29c455c1eeee58ccae90f30dff6a378d1c7bb0c013382722ba91

`define QX00 509'h809daccbda89f5414309d7471610e52f1ed06b37077baaba4f91c56a7a9f8b09c9c481da0183960a853bb53cc4384cdbf7d24ef9d54b5d4142930b33d7527e3
`define QX01 509'h1272fbdc27c1e8bb4bfa878616a86fb00cd1686b4ffeb70d1b4e4d2613e44b9664bc06f1f87ad9683a79bfb51d6803e3a841af5a0ec5bbaedb159619dfed5f1e
`define QX10 509'h25616e159857b6cedb6885b0a5a1bba132a05c35b97d21ec39bb61280948fc9335ff07d7efd8314ad31695ec387818498a28fe2914f24951525af24ece3d8f9
`define QX11 509'h11807e987a033cc404d5b7c44d74f0393c4568d6681387658e37165759e30f904e46b8f77905756c4d45f6d96fdb9f3ef18bbc89d58f1527f5dd9b5c76344f1a

`define TX00 509'h809daccbda89f5414309d7471610e52f1ed06b37077baaba4f91c56a7a9f8b09c9c481da0183960a853bb53cc4384cdbf7d24ef9d54b5d4142930b33d7527e3
`define TX01 509'h1272fbdc27c1e8bb4bfa878616a86fb00cd1686b4ffeb70d1b4e4d2613e44b9664bc06f1f87ad9683a79bfb51d6803e3a841af5a0ec5bbaedb159619dfed5f1e
`define TX10 509'h25616e159857b6cedb6885b0a5a1bba132a05c35b97d21ec39bb61280948fc9335ff07d7efd8314ad31695ec387818498a28fe2914f24951525af24ece3d8f9
`define TX11 509'h11807e987a033cc404d5b7c44d74f0393c4568d6681387658e37165759e30f904e46b8f77905756c4d45f6d96fdb9f3ef18bbc89d58f1527f5dd9b5c76344f1a

`define QY00 509'ha6a0618607608888346b865666940000dd661893d60628d12e071c3f05b3c52305f067a979439e074ae54a8871a1ad18589cde2331803ff6bd14dc517bb7d71
`define QY01 509'h15252e43e9615bc5a644517d36ccf9ac23c12f27049f9a4f6d78434162b037c1ba3d2f18092991d3afdffce38c606a37b8dd748ac5a782b49fb7f62d6a066991
`define QY10 509'hf5724b44eac77ea4498f6bb0a80cad03b67fa5338f016fc018f5065dec1d6ac89dd6cdad21a5f111ca210d14b197ac15b9b76dff0c987a913529a19628fac4d
`define QY11 509'h66edab04326e2a19fe1038c58811a5dbd446a69ee3ecb5749971217eecf5be14ba3f726dea8ae371083986f06b6fac9c973d0dbd6e6561249eeacd879d6f843

`define QY_00 509'haeb50e79ec3c21379a73a4f9357acf6bdb466c01fb81bff20098f3fefb55469320f7f44e48467105b1d07b7eaa0b90168d9ef253b758f01356bc3c8a104553a
`define QY_01 509'h3028bc15d86ed656a9a137c2f3f34aa7c999225878e43cc571bdc27d6058f9a83156a772ef0f1d1feb5f7ce55a699b3586487ca8e6104c01851b604eb9691a
`define QY_10 509'h5fe324bb08d52b1b854fbf9ef4022269022cdf624286790315ab09e014eba0ed89118e4a9fe41dfb3294b8f26a1591192c846277dc40b578dea77745630265e
`define QY_11 509'hee67c4fbc12e7fa5d0cef28a13fd2990e465ddf6ed9b334e952eeebf14134da16ca8e989d6ff2b9bf47c3f16b03d90924efec2b97a73cee574e64b53ee8da68

`define TY00 509'haeb50e79ec3c21379a73a4f9357acf6bdb466c01fb81bff20098f3fefb55469320f7f44e48467105b1d07b7eaa0b90168d9ef253b758f01356bc3c8a104553a
`define TY01 509'h3028bc15d86ed656a9a137c2f3f34aa7c999225878e43cc571bdc27d6058f9a83156a772ef0f1d1feb5f7ce55a699b3586487ca8e6104c01851b604eb9691a
`define TY10 509'h5fe324bb08d52b1b854fbf9ef4022269022cdf624286790315ab09e014eba0ed89118e4a9fe41dfb3294b8f26a1591192c846277dc40b578dea77745630265e
`define TY11 509'hee67c4fbc12e7fa5d0cef28a13fd2990e465ddf6ed9b334e952eeebf14134da16ca8e989d6ff2b9bf47c3f16b03d90924efec2b97a73cee574e64b53ee8da68

`define TZ00 509'haaaa90000c6356403120d4b063f1309347537b6a2e78173cd15fefc1fef6f449d917a4083e75f0f3034a39f8e452c2d119c42f891726cff5ec2ee7247402d55
`define TZ01 509'h0
`define TZ10 509'h0
`define TZ11 509'h0

