`define PX 1150'h249c309820e9d02ef25d7a834ab0b1400f72170f552fddf724f1fa92dac4a12f14edbbcd47be7689c17b3aa1f6f854df1a4c4fd6b6a4f653fc251820efcb13caf175caa79089a74e593f9d35ab8457de8654e9cce5d8064115ed248bd59a22e7665b033bb42b7be53b0932be73e84d468ef919e8e531d20a9dbfddaa494f77b68e6fcaada9376dec765544f791a28e1c
`define PX_ 1150'h15535a67df162fd10dae787e2d4f4ebff08e01242af0720ac97085712cf30629eb673d20bc64b826ad6a70010c98358603d6bbb8258b8fcaf5f755d11609e8b764457b8fbba0a3ac61402e15251c06ac7a830b8189a05e4b3717790d03bd3722ebb1ee59249e161c10ac55afb059590ed78d5ffe8acf6778324877b50405de6971a8f55260733cbe345595b319081c8f
`define PX3 1150'h33e506c862bd708cd70c7c88681213c02e562cfa7f6f49e380736fb488963c343e743a79d31834ecd58c0542e158743830c1e3f547be5cdd0252da70c98c3ede7ea619bf6572aaf0513f0c5631eca9109226c818420fae36f4c2d00aa7770eabe104181e43b8e1ae65660fcd3777417e4664d3d33f943c9d0937439f8e991103ab36a008f1fb9f1ab854f43c0a3cffa9
`define PY 1150'h1e20752166aa1a332f4176c073c9d091464c2f6dad85b654c01050e9a7d60445102ccda53f63bdd257abc9b65f3c386fc6146f07510daf67b1081028198302a55640511aea726d0e68196ab65940804919f402878f0146eeeaace089fbebc6928e4b50c297bc58c08f9517e8b0b74ac744ea545b142ce716a4cc1692a3c8c59b7b9a76fcfd490a93ba4988a86ece8ea8
`define PY_ 1150'h1bcf15de9955e5ccd0ca7c4104362f6eb9b3e8c5d29a99ad2e522f1a5fe1a313f0282b48c4bf70de1739e0eca45451f5580e9c878b22d6b741145dc9ec51f9dcff7af51c61b7ddec52666094775fde41e6e3f2c6e0771d9d6257bd0edd6b9377c3c1a0d2410d3940bc207085738a5b8e219c258c5bd4526c2b3c3ecca98c9084847e49030c61a016f06152023bdc1c03
`define QX0 1150'h9e28bba7f31cab72d845d67813f3f48929f6d2ee9ad9059c77ec33004fc794d0e9b607f53eac38e67c3840dea69627a71981ab03b287b485a69112ff7825cf35a4fdd10a9f09a1f2dad18c5340dc2968110421ddc71efd77574b52745904acf956ad348e13294c19b6b3f345b9521ead4f3fd72bb4e3d629b3a1eef0da7d329bc6e43f02afc0b2e4274dc1827db9339`define QX1 1150'h2c2231ef98bd991442ae70721c07fd84a97ecd3705973ec7f60ae6ca52163bd4e40ebdd1ed4060aa68f1e38ecf581164a896dcd3132c03ae5e95cd1e21e228e4ec9f5cbd1f10e845fea65c2dc1f8b53c260bc454706d51f6dc230c23d5e0a4a3adc8264dbf4f8624cbdd733f3816ec68c4d14e49b987afb3aa99d2f38ced63be8c3bf01ce14787912a4eebde3e20fe38`define QY0 1150'h1610a12736ffe208c1e957cb39b6867361204547cbc77d2ebf2f0dcebf40fb4f425b6a6b4a70d62cfe33df3d5f87a14695ed4bbea7303c71dbe42c5f6badbeb03a80a86153b3fd6395161c7a7a05d14b3f7c3f15a8f07eb30e61b36d482f265bb41a3e75ab9f126578fd647461d7a78469ca060310e05b207596b0c78f57f7e5ac473aab50ce487c264da20bad12e23e`define QY1 1150'h2d3fbb50dce34843c170bf636a43c393bd29435dd2c391f2deaa6d5b186b399b9e59590534bd6ec8ddf556fe2f6b25380b5fed5f74d9847f749494ad6bd3ad9b315c18b99e9d2e89d300ea624f075077c6c8e2a4190bc169728a1da3619e0ad4c394661c202ceed115266ab95c63d9a2035ae5f91b202d5d7e15e62471d2018408686e53d63765db2ca71bb6f5c36376`define QY_0 1150'h23dee9d8c9001df73e229b363e49798c9edfd2ebb458d2d32f3372354876ac09bdf98e82b9b2588370b1cb65a408e91e8835bfd0350049ad163841929a273dd21b3a9dd5f8764d972569aed0569a8d3fc15bb638c687e5d93ea2ea2b912833ae9df2b31f2d2a7f9bd2b823f9c269fed0fcbc73e45f20de625a71a497bdfd5e3a53d18554b8dc622e845d389efd97c86d`define QY_1 1150'hcafcfaf231cb7bc3e9b339e0dbc3c6c42d6d4d5ad5cbe0f0fb812a8ef4c6dbd61fb9fe8cf65bfe790f053a4d425652d12c31e2f6757019f7d87d9449a014ee7245f2d7dad8d1c70e77ee0e881990e133a0f12aa566ca322da7a7ff577b94f358e788b78b89ca330368f1db4c7ddccb3632b93ee54e10c2551f26f3adb83549bf7b051ac337344cf7e03bef3b4e74735`define TX0 1150'h9e28bba7f31cab72d845d67813f3f48929f6d2ee9ad9059c77ec33004fc794d0e9b607f53eac38e67c3840dea69627a71981ab03b287b485a69112ff7825cf35a4fdd10a9f09a1f2dad18c5340dc2968110421ddc71efd77574b52745904acf956ad348e13294c19b6b3f345b9521ead4f3fd72bb4e3d629b3a1eef0da7d329bc6e43f02afc0b2e4274dc1827db9339`define TX1 1150'h2c2231ef98bd991442ae70721c07fd84a97ecd3705973ec7f60ae6ca52163bd4e40ebdd1ed4060aa68f1e38ecf581164a896dcd3132c03ae5e95cd1e21e228e4ec9f5cbd1f10e845fea65c2dc1f8b53c260bc454706d51f6dc230c23d5e0a4a3adc8264dbf4f8624cbdd733f3816ec68c4d14e49b987afb3aa99d2f38ced63be8c3bf01ce14787912a4eebde3e20fe38`define TY0 1150'h23dee9d8c9001df73e229b363e49798c9edfd2ebb458d2d32f3372354876ac09bdf98e82b9b2588370b1cb65a408e91e8835bfd0350049ad163841929a273dd21b3a9dd5f8764d972569aed0569a8d3fc15bb638c687e5d93ea2ea2b912833ae9df2b31f2d2a7f9bd2b823f9c269fed0fcbc73e45f20de625a71a497bdfd5e3a53d18554b8dc622e845d389efd97c86d`define TY1 1150'hcafcfaf231cb7bc3e9b339e0dbc3c6c42d6d4d5ad5cbe0f0fb812a8ef4c6dbd61fb9fe8cf65bfe790f053a4d425652d12c31e2f6757019f7d87d9449a014ee7245f2d7dad8d1c70e77ee0e881990e133a0f12aa566ca322da7a7ff577b94f358e788b78b89ca330368f1db4c7ddccb3632b93ee54e10c2551f26f3adb83549bf7b051ac337344cf7e03bef3b4e74735`define TZ0 1150'h61074fffffffffffff40cfe87ffffffffffe7cc7fdfaffe119d7ffbf84858a6ffab0711fbdcd14f911a555cfc6f759ae1dcf47123cf79e10de3920dfa2b037daa44b9c8b3d5b505458034b52f5fa174ff280ab190879b73b2fb626726a8a5f5adf30e6b27366dfeb44a7791dbbe59aa997986188ffec67d2ff7aaa0b2aaa9dfffe73ffff65555555555255555555555`define TZ1 1150'h0