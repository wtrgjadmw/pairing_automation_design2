`define PX 440'h4d574b39e79d133d2aafc0a75a0221971b17b55511c7d5e0a2ff8ae5f14b3f6d8b5253c70104e0001f24bea4145e97a9e4aab2917857d
`define PX_ 440'hee2a8b502d7e98b881ddba686fb3b765cd1f59093a94d5b2d777f4af31e03da7125e86115997b7ccbc7c16c88a34f68d6109ff82e8252e
`define PX3 440'he805e1adb6d739b7800f41f60e0664c551471fff355781a1e8fea0b1d3e1be48a1f6fb55030ea0005d6e3bec3d1bc6fdae0017b469077
`define PY 440'h27993df832a7c852a07a287c8129756da32f0914d8608ec506ad9b386d8bedabbfd616e4d75c58f9f17842611ad599f869a128564da3ea
`define PY_ 440'hcb66c20b9950a199b40e8df6642a64119ba1cb49b350c44bdafa5225236903f22b3d9468f24bacd2ccf62051b0a5460f95b38255b206c1
`define QX0 440'h9d4e8568543ec797f9cb2f7f018effc1aa7a948a47b6c4de4eb8a319498e3cbfa590976f529aecdd8d0647031697260d22f4f99eea71a1`define QX1 440'h72bf4eae988fc592be7b4ea6e7e421f77d07d2aaeb5cb87151eab813b16b4783508c4138a09d0c7295c04c8f7f27384b0f8bfa72958a56`define QY0 440'h60a2d4e450c7e05d0cee221b0fd5210c62916eb913bce72f048959b0abd163d6f5f8b6a15e06be8e8f9c5befc91a977ad925d9f1f97d87`define QY1 440'h17e467c9fbf31555cab391c69eef3a07beeb98ec55763c6e27ba868f94cf2d62df4d8e41589a6c073175393fd0648e9496d26acacea589`define QY_0 440'h925d2b1f7b30898f479a9457d57eb872dc3f65a577f46be1dd1e93ace5238dc6f51af4ac6ba1473e2ed206c30260488d262ed0ba062d24`define QY_1 440'hdb1b9839d005549689d524ac46649f777fe53b72363b16a2b9ed66cdfc25c43b0bc61d0c710d99c58cf92972fb16517368823fe1310522`define TX0 440'h9d4e8568543ec797f9cb2f7f018effc1aa7a948a47b6c4de4eb8a319498e3cbfa590976f529aecdd8d0647031697260d22f4f99eea71a1`define TX1 440'h72bf4eae988fc592be7b4ea6e7e421f77d07d2aaeb5cb87151eab813b16b4783508c4138a09d0c7295c04c8f7f27384b0f8bfa72958a56`define TY0 440'h925d2b1f7b30898f479a9457d57eb872dc3f65a577f46be1dd1e93ace5238dc6f51af4ac6ba1473e2ed206c30260488d262ed0ba062d24`define TY1 440'hdb1b9839d005549689d524ac46649f777fe53b72363b16a2b9ed66cdfc25c43b0bc61d0c710d99c58cf92972fb16517368823fe1310522`define TZ0 440'hcfffffc34079613ab77498d1aac2680c12f2ba1744eacef1e5812a26f0b0e6214ec54b23657fa3341919d4d34851ff800ab5554005555`define TZ1 440'h0