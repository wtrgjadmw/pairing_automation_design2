`define PX 461'hb5d49be766a999724aaa974a7a442d5fc3360a30ad26a4c315f4d199d4585553689cb1e09a24daf9c216e6e09a1701858b10ad3abb628799ecc
`define PX_ 461'h9f80b86dee2c0be35ab2d1f6cef1ce772ead235affa3a2ee3253e290b9a7506e6364408a0ef07cf641e91b1f663e53cf1f99fd8544a82310bdf
`define PX3 461'hcc287f60df2727013aa25c9e25968c4857bef1065aa9a697f995c0a2ef095a386dd52337255938fd4244b2a1cdefaf3bf6875cf0321cec231b9
`define PY 461'h4130cee218a506410e633c3cd2ec04ea3892e58fcd50e6f8ff8380872796f8efb61b3406201569d05b56a6381fc1b1d37baa6d312627e98517
`define PY_ 461'h151424767334b54f19477357d7c073b884e59ff32aff53941b8507c221b863632d09f3f2a47140152fe4a979c7e593a3772f003eceda82c12594
`define QX0 461'hacba575538ced6ec7e17045a987b8be7be3d80fa519ede4e323ee4b9dbe708ed8f9c83c781e70844934e2d9f28d6be151ee21d41b26a1299636`define QX1 461'h6df4e42bf37fb0566ddbc5c8d5b19a188f347be8c3fe47b909c3a609242ae7a14ce0396aa82de79cf945e2305d60a71fdad7a773f0c729cd939`define QY0 461'h51e8eaec9f7d4c1e3a540cdc794ce38b548577e157a301a58189d96661bad3197c05c31127422b49f739cbd8553f22d67f81dc333e24ebd4a76`define QY1 461'h95b036ed6cb0de668952e79ebd688a5ed309b72c7ab1d81b28ef58c3f711483e488fc3f46e388414f03e1d87bb63185ec6d527f3cebb19afbc4`define QY_0 461'h1036c6968b55859376b095c64cfe9184b9d5db5aa5527460bc6bedac42c44d2a84ffb2f5981d32ca60cc63627ab16327e2b28ce8cc1e5bed6035`define QY_1 461'hbfa51d67e824c6ef1c0a81a28bcd71781ed9765f32186f961f595b6696ee5d8383712e763adcd3db13c1e47844f23cf5e3d582cc314f90faee7`define TX0 461'hacba575538ced6ec7e17045a987b8be7be3d80fa519ede4e323ee4b9dbe708ed8f9c83c781e70844934e2d9f28d6be151ee21d41b26a1299636`define TX1 461'h6df4e42bf37fb0566ddbc5c8d5b19a188f347be8c3fe47b909c3a609242ae7a14ce0396aa82de79cf945e2305d60a71fdad7a773f0c729cd939`define TY0 461'h1036c6968b55859376b095c64cfe9184b9d5db5aa5527460bc6bedac42c44d2a84ffb2f5981d32ca60cc63627ab16327e2b28ce8cc1e5bed6035`define TY1 461'hbfa51d67e824c6ef1c0a81a28bcd71781ed9765f32186f961f595b6696ee5d8383712e763adcd3db13c1e47844f23cf5e3d582cc314f90faee7`define TZ0 461'haaaaabaaab2a5aaa5aa296beb6ca04290e1cd2745335b84eb7b74bd572005a3e33ff0d9556eaa80ffbfffdffffaaaaab5555553ffff55555555`define TZ1 461'h0