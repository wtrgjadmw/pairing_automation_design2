`define PX 315'h1ca92fff0921082c6cb8dbb4002921d1be5608696f1c18f8b3fff3fe4fd147718c47a2e1fe7896
`define PX_ 315'h4a590d2b67db548a78a90b0357c358e0d037a12390afec7496ae5e6546e13bafe5bbb5c5e31876b
`define PY 315'h15146e010a9552973bc16371615c742ad9f0fe9f21e81915a9d906fa5f7759ecce051415c614ed1
`define PY_ 315'h370f322a4dd8127603b3354d366976d3122c030b05b994ee781556aacc66f63a307b1bde3ceb130
`define QX00 315'h22feab58cfdf3467f6bc5a83e34b0049459f223bd0d6fa49ac463ff7ae204ee50d04ff564b94336
`define QX01 315'h184cc36247e2f33d462b4e9229eaa05228a25c304c7248b276130b833ee6710f811ad2cb1214b65
`define QX10 315'hd29953c531a796991d473d2b9b7f0cee4d92eb2b80c61a7900aca2870fc4dbe7a12076399977f3
`define QX11 315'h3507b2daaca422228a0faeec45edd783226c3058b63edfb377c86d247ad702bae4f94b81d3711c9
`define QY00 315'h359c19b069be847b2687195144ebc7e521688144ed5b771659e5e7d6002e448581a71491c734241
`define QY01 315'ha5ec197010be045e51d69b0f31403c8b21e18dfdb5a3f542de267382216783c63d4951b70b5e06
`define QY10 315'h1a3164cb351201d554b22bbc853acdb7f895c7e1ee4b8089df298ba0c0ccdd17f65988f6a4bf102
`define QY11 315'h52caff12ffaf0bf3064b91ad2d5baba417c319f4a9003416d08d3e697a3d48c3c1e401f74e5487
`define QY_00 315'h1687867aeeaee09218ed7f6d52da2318cab480653a4636edc80875cf2bb00ba17cd91b623bcbdc0
`define QY_01 315'h41c4de94576184c75a572f0da4b1e73539fee8ca4c476eaff40bf66d09c7d7ea9aab9ad8924a1fb
`define QY_10 315'h31f23b60235b6337eac26d02128b1d45f38739c839562d7a42c4d2046b11730f0826a6fd5e40eff
`define QY_11 315'h46f6f03a2872744e0f0fdfa3c4f03043aaa0d00add11aac2b4e589be943a7b9ac261efd48e1ab7a
`define TX00 315'h22feab58cfdf3467f6bc5a83e34b0049459f223bd0d6fa49ac463ff7ae204ee50d04ff564b94336
`define TX01 315'h184cc36247e2f33d462b4e9229eaa05228a25c304c7248b276130b833ee6710f811ad2cb1214b65
`define TX10 315'hd29953c531a796991d473d2b9b7f0cee4d92eb2b80c61a7900aca2870fc4dbe7a12076399977f3
`define TX11 315'h3507b2daaca422228a0faeec45edd783226c3058b63edfb377c86d247ad702bae4f94b81d3711c9
`define TY00 315'h1687867aeeaee09218ed7f6d52da2318cab480653a4636edc80875cf2bb00ba17cd91b623bcbdc0
`define TY01 315'h41c4de94576184c75a572f0da4b1e73539fee8ca4c476eaff40bf66d09c7d7ea9aab9ad8924a1fb
`define TY10 315'h31f23b60235b6337eac26d02128b1d45f38739c839562d7a42c4d2046b11730f0826a6fd5e40eff
`define TY11 315'h46f6f03a2872744e0f0fdfa3c4f03043aaa0d00add11aac2b4e589be943a7b9ac261efd48e1ab7a
`define TZ00 315'h33dc5fd4a7929af2c08b6741683a150213e2fe55d85e51fbde11a25ad421afd9017fd00bfcfffff
`define TZ01 315'h0
`define TZ10 315'h0
`define TZ11 315'h0
