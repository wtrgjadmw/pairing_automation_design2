`define PX 317'hf51413257fea3fada43f18861510bee5390d4c513e44f4688f9e996a778f5ae8c93589303aa4fbe
`define PX_ 317'h10788f01761e532184bd41856a8c44ac3098d2170e2e5004df9504d8cabc9d000bdd5c35a00daed
`define PY 317'h6c5ce93755377160a9d2e482d91cb843d5d7809b84e02e3ea820f8888901a987b40be5d399aeb02
`define PY_ 317'h992fb8efa0d1216e7f297588a6804b4d93ce9dccc793162ec712a5bab94a4e612106ff924103fa9
`define QX00 317'h1300def2362dd93bebae729066aaa923f3bfe8782ae33a68080dbdb14ae3544fe68f4c99f61a969
`define QX01 317'h5e0770702f67d338788d55af7799f00ef34d55c176c2faa9efc3fd011637b617a70f214349da5f2
`define QX10 317'h28b472596bc81481cf6c0990e11d83cc87e1e1565fdf6f64694d4326475aa1e07afcce04989b3e4
`define QX11 317'h2f2759912bbb488ae951cbd1669e0e0be9f016ab171e57c4d0974bb4de56caac7978982e13a65f0
`define QY00 317'h56807b04098f4345aa72ed2d9cfef87e09d730232d08a34b79d26e75be8ff95322716f70a0860fa
`define QY01 317'h1970833cd8b56b5bbfea08928b3643c082ea756d112bf265829562674ab952e184aa7d3ed9b9520
`define QY10 317'heb58f264825348325de546580d6e2e34b55343906a9a2589ab5abbfc1e63cea0adbcb2cf6f86eeb
`define QY11 317'h2e2950a0209dd2953a4eb2979bdd4a743e07cdbb6979765430ca27870e0a7721d442d3ae64ee160
`define QY_00 317'haf0c2722ec794f897e896cdde29e0b135fceee451f6aa121f5612fcd83bbfe95b2a175f53a2c9b1
`define QY_01 317'hec1c1eea1d53277369125178f466bfd0e6bba8fb3b475207ec9e3bdbf792a5075068682700f958b
`define QY_10 317'h1a33afc273b54a9ccb1713b3722ed55cb452dad7e1d91ee3c3d8e24723e82948275632966b2bbc0
`define QY_11 317'hd7635186d56ac039eeada773e3bfb91d2b9e50ace2f9ce193e6976bc344180c700d011b775c494b
`define TX00 317'h1300def2362dd93bebae729066aaa923f3bfe8782ae33a68080dbdb14ae3544fe68f4c99f61a969
`define TX01 317'h5e0770702f67d338788d55af7799f00ef34d55c176c2faa9efc3fd011637b617a70f214349da5f2
`define TX10 317'h28b472596bc81481cf6c0990e11d83cc87e1e1565fdf6f64694d4326475aa1e07afcce04989b3e4
`define TX11 317'h2f2759912bbb488ae951cbd1669e0e0be9f016ab171e57c4d0974bb4de56caac7978982e13a65f0
`define TY00 317'h56807b04098f4345aa72ed2d9cfef87e09d730232d08a34b79d26e75be8ff95322716f70a0860fa
`define TY01 317'h1970833cd8b56b5bbfea08928b3643c082ea756d112bf265829562674ab952e184aa7d3ed9b9520
`define TY10 317'heb58f264825348325de546580d6e2e34b55343906a9a2589ab5abbfc1e63cea0adbcb2cf6f86eeb
`define TY11 317'h2e2950a0209dd2953a4eb2979bdd4a743e07cdbb6979765430ca27870e0a7721d442d3ae64ee160
`define TZ00 317'hfa735dd909f76d30d703a5f48062fc6e9659e197b38cbb9290cc61bcbdb408172aed1a9a254d555
`define TZ01 317'h0
`define TZ10 317'h0
`define TZ11 317'h0
