`define PX 318'h2c4f942191b5adf67c4fd50f1a56827dccffb1b3b0baef315e3fb866f05b20489112a95b4723e2bf
`define PX_ 318'h7151979f57ed769e780e36088f4f0b23c676eb25662b92be7fff35ebdfbf766f424ca4693177ec
`define PY 318'h128b4a3cdf573bbe6e7fd29e943baa12439cff1c38673048d8f6cfb103911a5e3b51680b6ae83075
`define PY_ 318'h1a359b7c51b65faeac4810a68eaa2776ad2929829db9ea7b43c8e7ebd8a9c560c5038df4456d2a36
`define QX00 318'h2924322cfc9c9476823c9939fd64afcba73c3e2a2160f0cd9f36043ea62146fac4f6509cffff3aaa
`define QX01 318'h231b5db64e977f624dc8fb3014088d1b1b8e651601ce3615c47188e745b9539ac9e04d39704955c5
`define QX10 318'h221003670cdec5d4043974c8bb6ce113fc0ce94dd47d30003c2f9a20f63d440476b09d18c405ce79
`define QX11 318'h231b42544f477e4e21181a4a9b4988442391affc469d97c5189dbe2878533f1fb48e7f88a327c993
`define QY00 318'h25a134b7879fc3e73f21ca438ebecfec149583831c1a9b58458e072eb28c6cd59d0df4cc79b65933
`define QY01 318'habc923162d7293bf55450fc9f5ed84ebd5db2d8f54b584378844527eb7b37721f6d78e067b9a2cc
`define QY10 318'h1e7cc2236bc917f7fdaf606258680f3c2bb17d53a0bb27fe9d04d9bcc42854de217707d2393d444f
`define QY11 318'h7e53f41e456b66f4daf22ef930406e69b3990c90eb1ef2b9359ae119a571e861a0888761a2d59
`define QY_00 318'h71fb101a96dd785dba619019427019cdc30a51bba067f6bd731b06e29ae72e963470133369f0178
`define QY_01 318'h22045387ce367231257392488386f93a336875c5e0d5c280a43b7274f0bfa84ce0e77d1f489bb7df
`define QY_10 318'he442395c54483751d1882e2ca7dc24cc514ab4b3565f2c57fbadde018128ae0deddee2d7718165c
`define QY_11 318'h2cb90079ef2944b6ab7a34223352cd820a2aef0e0d1268d4f12c5deecaa088a07a3aed773a3b2d52
`define TX00 318'h2924322cfc9c9476823c9939fd64afcba73c3e2a2160f0cd9f36043ea62146fac4f6509cffff3aaa
`define TX01 318'h231b5db64e977f624dc8fb3014088d1b1b8e651601ce3615c47188e745b9539ac9e04d39704955c5
`define TX10 318'h221003670cdec5d4043974c8bb6ce113fc0ce94dd47d30003c2f9a20f63d440476b09d18c405ce79
`define TX11 318'h231b42544f477e4e21181a4a9b4988442391affc469d97c5189dbe2878533f1fb48e7f88a327c993
`define TY00 318'h71fb101a96dd785dba619019427019cdc30a51bba067f6bd731b06e29ae72e963470133369f0178
`define TY01 318'h22045387ce367231257392488386f93a336875c5e0d5c280a43b7274f0bfa84ce0e77d1f489bb7df
`define TY10 318'he442395c54483751d1882e2ca7dc24cc514ab4b3565f2c57fbadde018128ae0deddee2d7718165c
`define TY11 318'h2cb90079ef2944b6ab7a34223352cd820a2aef0e0d1268d4f12c5deecaa088a07a3aed773a3b2d52
`define TZ00 318'h133f1a46cef26492e5381cbadd1a2e770f39d76129dee53be340486323c52040ffab0a004faaa555
`define TZ01 318'h0
`define TZ10 318'h0
`define TZ11 318'h0
