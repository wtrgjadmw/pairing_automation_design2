`define PX 1032'h25f400f1f53d085114ae9500a4a2ad82816ca62943f92df576453fc0755247bf6fd7a709d913979bc17ec0faf91a7e32b676a567e58c2ca132f3778edc9c603dc2ba159b519a176503b662a2580e3ad7085e8194f628336530bba44d0812034712b711924e7dbc74e25150e5c2bf02d413c582e9d05bf25c5277efab7591e765b
`define PX_ 1032'hc44f61456f52b1cf9fc81d0ea81b354b87b60e90756302daf8a2a2b7140cd4fa7576d6453a6c23368d4e16184411dc85c7e84d9b334819fb8de6935b644a245f9e598c91ab5854604027ae54a53698c9c4da713bcef147c934744b20907ee22b8eb7397185bd79af073040404e7d0fd3141927d132fa40da402dd7aff3518c3450
`define PY 1032'h4f0075a5b4466cf30f68de71a7c400005be0e7b9663871a2bc2ac93494341f0a1810b3ca70010d8e6d14369167b4719cb9a455b8da246f9d240c8a800c1475e5e5670b2dbff34dd7c0de93b49bd8ef35c815698638f23d4d4af6b264bf8556960e3b80d1e9bb5958e0de8df1d8e3d2be6c211de828fbb4ccc6c0baaa070a7b2835
`define PY_ 1032'h77ae2baeda601561a1aa27ed0aa1602353ebf139a36a241793dc2d7e872dda6c54639ceb67fc4f21dc51cb968bef12cc39ab6238d77c6d287d09405445ff747d951e22bda07ea7fecf8480ca2ede8d416d4aefcee5618db23c895300a17aabc9f1a729b8c0e9fc1d7476c75cd1c52d41e9346217a7044b333e949c00a3a02f8276
`define QX00 1032'hc5b29031647944f1ab30cbbe1f90b8d19679df9f3aa0b1b01c54402f73bfc427e554c00b88985759cd3a570cf9b4c0e96456907853af28cc694e662f6c7d1743a91dc143d006366cbe3bb7b5f956d8ffa204fb8aafc5e7a7e3e9d45f1acd70d5546c01d7f20d0458d383f40c05d75bb4e32fa52f616d77a52c046fa6fd015bde5b
`define QX01 1032'h8b39fe89131840e678bd8dca36e7da289d18e3d8cc29aebe230f083f3b925246d2a1fc5fd7ed2bfc2233e5317354e33a360265803e34e11030908c88e8ad8cc4f5f90b02c79c28b4bd69bd5648501bceda058435c051ffc94da127860c4b63ff627125e1a1eefc3fc3361b7da6ddd6bdd9dabe2e1aef63c4a530ed29d411a858ac
`define QX10 1032'hb333dd2fd759922575819772e6681b348fd10f0eba68004b4400e4419a35296e98e3de565be5a1425222a44c14f5ad92d01f283f1cc4cbcf32da797eea333a46e0e879cf7b2cf94b9276b1bfdf57b9b32d96bc3e32756fdca87a1c0ad10945c7df7ca4919d5119a3792f1e12fd86bb44711510b735925819fbdf0b827a748b0f4f
`define QX11 1032'h58205f7cc572acd04916dbd0d1b42cf1bd1cc1688454a3233d79b7ad3851d2b66948d2a7751c07988a58a6571467a05dd4a73c8ec8c31b70a8762897ee0f0365e75c8eea78705c3ebed29523354c7666425025e404ef570ea3769058ca780685bb8ba21643b158635ff25c2f2bb4b72e22af6508981421fe6b36dead3becf59fa7
`define QY00 1032'hc0eacac68f644195553072adcbc31e28917c34b1ee14e227be818c64f154f0e1f87881689edfcd471c51ee4f2bb596f012a189eeb7ad7ffc2ba06a598328fee4b3c2525083150ecfcbb1c092019224700c0dfbc63ef70d78635f95c629fb0c65a41c2e485d010195b563d651eec2b18ca5cc9bcc9151a22ff7f542b2cfaa51bdc0
`define QY01 1032'h54e2d8b03204be64d22350ae0dbf494ac35145234eb82b7ea36548a3bdd234a275e4c2d9eb1104d1535b3be23f454c21e23d4bac6844e93b03a32e22cf6168448a7386a659daa9586e7684033ca43811a5da7bfba3554ce46891157bc92f6d6e4f471192d19f53189cb25fe8e1488d4a51efdd2e923c77739ef3a6d27471b4311d
`define QY10 1032'h5d6936afef36f22bcc5def4b52b11a4ca9f61f95cb8d70410a88dc56d4bc760b909bed60c8c1c0702dd3e856c239bbe29bc459d8170743f8d8217711c9023f6e27b53a4f940e30137b49a764a869f25406350ee0523fe4b8b976bcc76d3edbd39c795ca665ac9ad3ea678bf8ec4f8f1463122c82ecdace254bc05eb020fbee7664
`define QY11 1032'h68cb4be456c22036ca553de0e8d4191852c628daa9339a8e7a862fffce682f02d255928d8303b155b65312c208a6c4092c660612a4c6da29f062cd9e1d71eb0ac6b619d797b6819e0d3c805bfa21902ccb7823707c3297f7882d8660b5ce59b9d2505f3a64e7361eee352e6df630d38dd2c3e149944ffd548d8c3ee0dbecaa61e1
`define QY_00 1032'h5c3d68dff4240bf5be293b0e6a241fb1e50a4411b8db39291856a4e2a0d089473fbcf4d391d8f692d1413d8c7eded78e0ae2e02f9f35cc97575607aceeaeb7ec6c2db9add5ce706c4b153ecc925580729525d8edf5cbd8724206f9f3704f5fa5bc67c424da453e09ff17efcbbe64e73af88e4333eae5dd00d6013f7db0058eceb
`define QY_01 1032'h71cbc8a45ca1c3efdeefb5b0a4a616d8ec7b93cfbaea6a3baca1ae0f5d8fc4d3f68f8ddbecec57def60ac645b45e384711126c45495bf38a9d729cb182b2821ef011a74506974c7e21ec907b8e1344658f85dd597afe7e1b1eeeefe997d094f1b09b98f7d906025db8a2f565c96072b60365a2d13dc3888c6661afd83638f6798e
`define QY_10 1032'h69456aa49f6f9028e4b517135fb445d705d6b95d3e152579457e1a5c46a5836adbd863550f3b9c401b9219d13169c886578b5e199a9998ccc8f453c28911aaf552cff39bcc63c5c315196d1a224d8a232f2b4a74cc13e646ce09489df3c1268c63694de444f8baa26aedc955be5970ebf243537ce32531dab994f7fa89aebc3447
`define QY_11 1032'h5de3557037e4621de6bdc87dc991470b5d06b018606efb2bd580c6b34cf9ca739a1ebe2854f9ab5a9312ef65eafcc05fc6e9b1df0cda029bb0b2fd3634a1ff58b3cf1413c8bb743883269422d095ec4a69e835e4a2213307ff527f04ab31a8a62d924b5045be1f57672026e0b4782c7282919eb63bb002ab77c917c9cebe0048ca
`define TX00 1032'hc5b29031647944f1ab30cbbe1f90b8d19679df9f3aa0b1b01c54402f73bfc427e554c00b88985759cd3a570cf9b4c0e96456907853af28cc694e662f6c7d1743a91dc143d006366cbe3bb7b5f956d8ffa204fb8aafc5e7a7e3e9d45f1acd70d5546c01d7f20d0458d383f40c05d75bb4e32fa52f616d77a52c046fa6fd015bde5b
`define TX01 1032'h8b39fe89131840e678bd8dca36e7da289d18e3d8cc29aebe230f083f3b925246d2a1fc5fd7ed2bfc2233e5317354e33a360265803e34e11030908c88e8ad8cc4f5f90b02c79c28b4bd69bd5648501bceda058435c051ffc94da127860c4b63ff627125e1a1eefc3fc3361b7da6ddd6bdd9dabe2e1aef63c4a530ed29d411a858ac
`define TX10 1032'hb333dd2fd759922575819772e6681b348fd10f0eba68004b4400e4419a35296e98e3de565be5a1425222a44c14f5ad92d01f283f1cc4cbcf32da797eea333a46e0e879cf7b2cf94b9276b1bfdf57b9b32d96bc3e32756fdca87a1c0ad10945c7df7ca4919d5119a3792f1e12fd86bb44711510b735925819fbdf0b827a748b0f4f
`define TX11 1032'h58205f7cc572acd04916dbd0d1b42cf1bd1cc1688454a3233d79b7ad3851d2b66948d2a7751c07988a58a6571467a05dd4a73c8ec8c31b70a8762897ee0f0365e75c8eea78705c3ebed29523354c7666425025e404ef570ea3769058ca780685bb8ba21643b158635ff25c2f2bb4b72e22af6508981421fe6b36dead3becf59fa7
`define TY00 1032'h5c3d68dff4240bf5be293b0e6a241fb1e50a4411b8db39291856a4e2a0d089473fbcf4d391d8f692d1413d8c7eded78e0ae2e02f9f35cc97575607aceeaeb7ec6c2db9add5ce706c4b153ecc925580729525d8edf5cbd8724206f9f3704f5fa5bc67c424da453e09ff17efcbbe64e73af88e4333eae5dd00d6013f7db0058eceb
`define TY01 1032'h71cbc8a45ca1c3efdeefb5b0a4a616d8ec7b93cfbaea6a3baca1ae0f5d8fc4d3f68f8ddbecec57def60ac645b45e384711126c45495bf38a9d729cb182b2821ef011a74506974c7e21ec907b8e1344658f85dd597afe7e1b1eeeefe997d094f1b09b98f7d906025db8a2f565c96072b60365a2d13dc3888c6661afd83638f6798e
`define TY10 1032'h69456aa49f6f9028e4b517135fb445d705d6b95d3e152579457e1a5c46a5836adbd863550f3b9c401b9219d13169c886578b5e199a9998ccc8f453c28911aaf552cff39bcc63c5c315196d1a224d8a232f2b4a74cc13e646ce09489df3c1268c63694de444f8baa26aedc955be5970ebf243537ce32531dab994f7fa89aebc3447
`define TY11 1032'h5de3557037e4621de6bdc87dc991470b5d06b018606efb2bd580c6b34cf9ca739a1ebe2854f9ab5a9312ef65eafcc05fc6e9b1df0cda029bb0b2fd3634a1ff58b3cf1413c8bb743883269422d095ec4a69e835e4a2213307ff527f04ab31a8a62d924b5045be1f57672026e0b4782c7282919eb63bb002ab77c917c9cebe0048ca
`define TZ00 1032'h39515eab71597dab4eecf9a14d9a9fdc5033270cf65d6a45aff9094ce49e0689938baf4a2802a34fb699fdd80c5c7b970cb0480e4e5f233a5eea352badec159c857ad2149f8e0a296f9ceb8135488388ca9fa6aae1ac3500787ffa9a9efffda0001d5575555aaa89aaaaaab15556ffffaaaa80002ffffffffaaaa9555555555555
`define TZ01 1032'h0
`define TZ10 1032'h0
`define TZ11 1032'h0
