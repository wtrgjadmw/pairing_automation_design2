`define PX 559'h28a6152fcde32c9c440da0a0891fae4717a41b77440ca8de328004baf446e79ca96f276c668e9a8a22a370741c6fabe9e7b384b00842a8f123e77b9da10891d48991f2bab402
`define PX_ 559'h2cc9ee90821b5d3f0de1e624e0015ad704ceb671df8b2b400542511250a908b51a2080a740072b4b51eecb7ac6e401b7285686afa9ce7136595117c5367739839656c24651e9
`define PY 559'h447d75c6263da87d6e1ad7f2c39356ac1aef0c0ad3a0fe4654ee37b3d3a0b04219ee705dc1ea7f0617e84e23ccdecdaa1f0e253c41430713f9c0ed47fc4217e6c20596f229b2
`define PY_ 559'h10f28dfa29c0e15de3d4aed2a58db2720183c5de4ff6d5d7e2d41e19714f400fa9a137b5e4ab46cf5ca9edcb1674dff6f0fbe62370ce13138377a61adb3db3715de31e0edc39
`define QX00 559'h4965e279fcee4078339730e793926831070bf39fe877b098230a873872e98ba9a2bd7fc8ddd0e0b71b5d331861a745e8167dc4d10fc72307597644a45ca62ec48e3bdeb57cd9
`define QX01 559'h21e92a2e3fa5b458d21480b5e013d1858e25cc1e8d4503ff25a62cd67a454d49bf77719440edb7c20967e4c56c1018b672e3cc594e8ce0156e4dc03d02d3d32f699d7dae226d
`define QX10 559'h24cad2fdf6663f87aa89e10e9eb85a37c5f4b7f55c43774bb60a20d301e7aa9309cc48fc709bb7660457d210da45463ac2b617ea351fd0cc1d6d85dff73ffaf754801b3163c0
`define QX11 559'h21f505f984e0264236d1f1d6be0ded73b03b9a9bdfd6f40641f41a33897f516ffe1e4e2078ff24a52b097964b225bc843043f8054f5089cec709e04f02458c095e422130570f
`define QY00 559'h4861b77fa2c9e281e2599b22fc7b854869628ce478e9f08974ebdff8f65602d0f719d2e8eb85ce2a55608d74a1a065ffd392272121b18e492567f7ad04c23df5c4cbf34b6f0b
`define QY01 559'h1e03f42705c5b1a2c0a2c17d3788a00be294d32c617889e646bb3cc43cb8965d19d2baa23c48b05ec0684e7340aa1bbdd1d86b3e18e1bb4103b1e0de58e37d169d55605a44e7
`define QY10 559'h4706b3b7908015b7308b4a2d53510fa9372b9f704822207a9f71ebbd47662078a5dbc20917f71487eb354a7cbd449be46df38a9e49086a135f5aa0d7cda0f455a818d82ddd28
`define QY11 559'h3078e7ca8adaac7d32a5cae22a511ee03329715f2ce0bc9abacd8e72969e24c2eccd0c0020039b87d471abc6429e52ea8a09f110ac85b934353fc8d1f90aa9a1674f2f287b80
`define QY_00 559'hd0e4c40ad34a7596f95eba26ca583d5b3104504aaade394c2d675d44e99ed80cc75d52abb0ff7ab1f31ae7a41b347a13c77e43e905f8bde57d09bb5d2bd8d625b1cc1b596e0
`define QY_01 559'h376c0f994a38d838914cc5483198691239ddfebcc21f4a37f1071909083759f4a9bced716a4d1576b429ed7ba2a991e33e31a021992f5ee67986b2847e9c4e41829354a6c104
`define QY_10 559'he695008bf7e742421643c9815cff974e5473278db75b3a398506a0ffd89cfd91db3e60a8e9eb14d895cf172260f11bca21680c16908b0141dddf28b09ded70277cfdcd328c3
`define QY_11 559'h24f71bf5c523dd5e1f49bbe33ecfea3de9496089f6b717837cf4c75aae51cb8ed6c29c1386922a4da0209028a0b55ab686001a4f058b60f347f8ca90de7521b6b89985d88a6b
`define TX00 559'h4965e279fcee4078339730e793926831070bf39fe877b098230a873872e98ba9a2bd7fc8ddd0e0b71b5d331861a745e8167dc4d10fc72307597644a45ca62ec48e3bdeb57cd9
`define TX01 559'h21e92a2e3fa5b458d21480b5e013d1858e25cc1e8d4503ff25a62cd67a454d49bf77719440edb7c20967e4c56c1018b672e3cc594e8ce0156e4dc03d02d3d32f699d7dae226d
`define TX10 559'h24cad2fdf6663f87aa89e10e9eb85a37c5f4b7f55c43774bb60a20d301e7aa9309cc48fc709bb7660457d210da45463ac2b617ea351fd0cc1d6d85dff73ffaf754801b3163c0
`define TX11 559'h21f505f984e0264236d1f1d6be0ded73b03b9a9bdfd6f40641f41a33897f516ffe1e4e2078ff24a52b097964b225bc843043f8054f5089cec709e04f02458c095e422130570f
`define TY00 559'hd0e4c40ad34a7596f95eba26ca583d5b3104504aaade394c2d675d44e99ed80cc75d52abb0ff7ab1f31ae7a41b347a13c77e43e905f8bde57d09bb5d2bd8d625b1cc1b596e0
`define TY01 559'h376c0f994a38d838914cc5483198691239ddfebcc21f4a37f1071909083759f4a9bced716a4d1576b429ed7ba2a991e33e31a021992f5ee67986b2847e9c4e41829354a6c104
`define TY10 559'he695008bf7e742421643c9815cff974e5473278db75b3a398506a0ffd89cfd91db3e60a8e9eb14d895cf172260f11bca21680c16908b0141dddf28b09ded70277cfdcd328c3
`define TY11 559'h24f71bf5c523dd5e1f49bbe33ecfea3de9496089f6b717837cf4c75aae51cb8ed6c29c1386922a4da0209028a0b55ab686001a4f058b60f347f8ca90de7521b6b89985d88a6b
`define TZ00 559'h2a8ffc3fb0017624ae10793a96def6e1e38d2e16dc682be1c83daa32bb100fae3c7057ec596a3a2a8b6dc4111cac525eeff5f4a04deee5d882c76c9d288034a7e0174afefa15
`define TZ01 559'h0
`define TZ10 559'h0
`define TZ11 559'h0
