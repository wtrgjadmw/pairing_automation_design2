`define PX 446'h23f29a3ddc00a4b60b8dab725e752b8027442e426c263313033c610ee3118748ba5eaa2001034e453ce74dbd869df7cba82224707073b3c7
`define PX_ 446'h18ec46bd4cc5407f148217d70735aabfd95176751ddccb1f0c39453cd7b58eb9c7efc3a3e1377fa91a06f76b3ed5be0088f9dbb63a3cf6e4
`define PX3 446'h2ef8edbe6b3c08ed02993f0db5b4ac407536e60fba6f9b06fa3f7ce0ee6d7fd7accd909c20cf1ce15fc7a40fce663196c74a6d2aa6aa70aa
`define PY 446'h11cf7b046fe41c150fa7607243eed9044605cf5314391d3f7dabb4073a99600c4dca0a0312059b43b304c11d7266d645868147503a1e2956
`define PY_ 446'h2b0f65f6b8e1c920106862d721bbfd3bba8fd56475c9e0f291c9f244802db5f6348463c0d03532aaa3e9840b530cdf86aa9ab8d670928155
`define QX0 446'h2833f24971f57d09d759864ae026f766d787a7d467e5b5823a8b49f0675ca23fb665147c60866b400b5f3a06daab0b85e477017b00fcdf99`define QX1 446'hf9116e6a02660d134162fe2adfc3e4ce83c346d0da55c0f747373e1c1c7c37a3fd3256916c607537789152750a03adb3b61fcc0e88aa3db`define QY0 446'h24c894f18bc44d729e5f59523b62149fad1c14b3e510628ef05fc6362f7fe9f9aa0310d1b2b2724984ff30e52736de1f448fa2afafc1498`define QY1 446'hece8ac5182d2081221d8c0e2f2e57e19ced5ffb6a7d33b54eecdd4717a69102e366691526836126e6257c8f3d88ce37735d086fa3a250ec`define QY_0 446'h3a9257ac1009a05df629cdb441f4b4f605c3e36c4bb1f809206fa9e857cf1762e7ae3cb6c70fa6c9be9e521a730047ea3cd305fbafb49613`define QY_1 446'h2e1056361098c4b3fdf2373b367c7e5e63a844bc1f85ca7cc088c904a32084ff9ee804aebbb76cc770c8c89987eae794bdbef7b7070e59bf`define TX0 446'h2833f24971f57d09d759864ae026f766d787a7d467e5b5823a8b49f0675ca23fb665147c60866b400b5f3a06daab0b85e477017b00fcdf99`define TX1 446'hf9116e6a02660d134162fe2adfc3e4ce83c346d0da55c0f747373e1c1c7c37a3fd3256916c607537789152750a03adb3b61fcc0e88aa3db`define TY0 446'h3a9257ac1009a05df629cdb441f4b4f605c3e36c4bb1f809206fa9e857cf1762e7ae3cb6c70fa6c9be9e521a730047ea3cd305fbafb49613`define TY1 446'h2e1056361098c4b3fdf2373b367c7e5e63a844bc1f85ca7cc088c904a32084ff9ee804aebbb76cc770c8c89987eae794bdbef7b7070e59bf`define TZ0 446'h3211f04d73a1acadff03cb69a5529bfff6a5b4875fd01cdf08a59b44538e9fd7db1923c1dc53211a911bad73a8c4a33cee3ffd9554f5555`define TZ1 446'h0