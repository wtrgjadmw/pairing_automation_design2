`define PX 559'h21a7d414d9f2d0f7435b751e365dbbcbc46e4f7b7cdc3e5993f6f99c9daed394af0397d91373889ea31909b0c1b46ff28beaca232469c684c5b0a53d2bd101a0bcfee4ee6444
`define PX_ 559'h33c82fab760bb8e40e9411a732c34d525804826da6bb95c4a3cb5c30a7411cbd148c103a93223d36d179323e219f3dae841f413c8da753a2b787ee25abaec9b762e9d012a1a7
`define PY 559'h7063b4b9fd306eb4b40c85573878342b7944316e022b7b1ec0e59d456cebf1b4e7906e12fd87ada579a1e760b8a4388e76a8bf6baab0545f4035653732d275fb9fb2045b520
`define PY_ 559'h4e69c874b02b82f006aebe6ff59985db64de8ed243751c6c4bb3fbf8ee2131367516a13276bd4afb1cf81d78d7c96a18289f7f68f76614e189353d0f6452a3f865ed94bb50cb
`define QX00 559'h3b38b38392df8f9f40276735bd2e4d3eafa163e5d251fdb855c8b0e538cc261952b353996f74789fd1ffe81c432162d312d0ff07b0fc449f87df205ff509219ba05d5897c800
`define QX01 559'h3e9e4bdc5eac811734b276474f4dbba02b694232a1ff31dea51d1b3bd740eaf5a00fba73e7529a4938e9a80e65b2dc42f876f7af4a7c0f97beb67192ba514152e21fa63180c6
`define QX10 559'h3bef499a1b3aa2f46e546deca20b12093cdf614e31f172dcf60c7cfed1f8e80c322b2afcd1bbbba598066e06d6c773931bfb80bf0dbf6550eba3b693f5c13c391805037063b3
`define QX11 559'h387ae000c3831b66dfdf9838060daa248a674862806e7e217cae4d465c112fcc9d2617903ca9fff44a8ad237fc9417ee8d86513d6be025e42a6cebe7558ca65042b4bba6db34
`define QY00 559'h19d6ddca464333f6ce663e6d1b3bc8d0900abdaba847b3cd7aefd4ca693dcf34978a2da6d8ca82e7692fb68843476bc6af25684fe2118b80eba9989f91e75cd1fe2cd1dfc294
`define QY01 559'hb86f51cd00c1c1ab232f3df8d316bb0df5a16d052bf16d565df064df36120f7e33d5f37b8f48b1a625bb15faff89cfd63615de6bca77f6c8b8200ba2b892a5a182088aa4052
`define QY10 559'h1bd2dcda8f6a68ad5d2c1b47e8b2175f442d59c83fa18a40c96b9599df8554c9df8af74d2e52e1277033b5961e3028b2a73421f952e5fb66180a38ab8041f9bfc2f56904ee93
`define QY11 559'h32e46a106ba984710151042250fed6ab01d354b596ac2e224017a7fb4bae8a335e0c243c260c4b6e3a990fd011fc4fbf626c5eb49d2f3abe15dbb3ca4740d41b129c8ab579a7
`define QY_00 559'h3b9925f609bb55e4838948584de5404d8c68143d7b502050bcd28102dbb2211d2c057a6ccdcb42ee0b628566a00c41da60e4a30fcfff8ea6918efac345986e8621bbe3214357
`define QY_01 559'h49e90ea37ff26dc09fbc92e5dbef9d6d3d18bb18d0d8bd48d1e34f7f518ecf59e05248dbeda13abb12368a8f335b10a3aca8ad78f5699abaf1b692a8abf6a0fe07c82c56c599
`define QY_10 559'h399d26e5c094212df4c36b7d806ef1bed8457820e3f649dd6e56c033656a9b87e404b0c67842e4ae045e8658c52384ee68d5e9665f2b1ec1652e5ab7573dd1985cf34bfc1758
`define QY_11 559'h228b99afe455056a509e82a3182232731a9f7d338ceba5fbf7aaadd1f941661e658383d780897a6739f92c1ed1575de1ad9dacab14e1df69675cdf98903ef73d0d4c2a4b8c44
`define TX00 559'h3b38b38392df8f9f40276735bd2e4d3eafa163e5d251fdb855c8b0e538cc261952b353996f74789fd1ffe81c432162d312d0ff07b0fc449f87df205ff509219ba05d5897c800
`define TX01 559'h3e9e4bdc5eac811734b276474f4dbba02b694232a1ff31dea51d1b3bd740eaf5a00fba73e7529a4938e9a80e65b2dc42f876f7af4a7c0f97beb67192ba514152e21fa63180c6
`define TX10 559'h3bef499a1b3aa2f46e546deca20b12093cdf614e31f172dcf60c7cfed1f8e80c322b2afcd1bbbba598066e06d6c773931bfb80bf0dbf6550eba3b693f5c13c391805037063b3
`define TX11 559'h387ae000c3831b66dfdf9838060daa248a674862806e7e217cae4d465c112fcc9d2617903ca9fff44a8ad237fc9417ee8d86513d6be025e42a6cebe7558ca65042b4bba6db34
`define TY00 559'h3b9925f609bb55e4838948584de5404d8c68143d7b502050bcd28102dbb2211d2c057a6ccdcb42ee0b628566a00c41da60e4a30fcfff8ea6918efac345986e8621bbe3214357
`define TY01 559'h49e90ea37ff26dc09fbc92e5dbef9d6d3d18bb18d0d8bd48d1e34f7f518ecf59e05248dbeda13abb12368a8f335b10a3aca8ad78f5699abaf1b692a8abf6a0fe07c82c56c599
`define TY10 559'h399d26e5c094212df4c36b7d806ef1bed8457820e3f649dd6e56c033656a9b87e404b0c67842e4ae045e8658c52384ee68d5e9665f2b1ec1652e5ab7573dd1985cf34bfc1758
`define TY11 559'h228b99afe455056a509e82a3182232731a9f7d338ceba5fbf7aaadd1f941661e658383d780897a6739f92c1ed1575de1ad9dacab14e1df69675cdf98903ef73d0d4c2a4b8c44
`define TZ00 559'h2a8ffc3fb0017624ae10793a96def6e1e38d2e16dc682be1c83daa32bb100fae3c7057ec596a3a2a8b6dc4111cac525eeff5f4a04deee5d882c76c9d288034a7e0174afefa15
`define TZ01 559'h0
`define TZ10 559'h0
`define TZ11 559'h0
