`define PX 381'hdf6a6a7f6b9ba536f9a25e48ef939a0f0fe50fd2f36db4d973a84e5a2fd43a3fd6c794b8a7e85ef6ef01754fb3ea12a
`define PX_ 381'hc0a6b4242c62c46db8181d1b45273367378fa87c44e3771cff64dbb53b3b280213f86b326d57a104b0ee8ab04c10981
`define PX3 381'hfe2e20daaad486003b2c9f769a0000b6e83a7729a1f7f295e7ebc0ff246d4c7d9996be3ee2791ce92d145fef1bc38d3
`define PY 381'h11504983887e59d4acc852e905b3b9ac7f42445389accba3393d6cdb12684fe3c9adfebf59dfc92b71ba8c62cfe1d613
`define PY_ 381'h8b0c866b1018cc59e5354cd3d97f32ae535073169d8471c2df365c5e448a64054fe013f577436d44844739d301dd498
`define QX0 381'h10b8501b92fe9329d24e30191ee6b5d10034a5eedfa61f71daaa1975e1b40b7c91a33c5021eff7f29fe39f429fa0a269`define QX1 381'h4ec8b6dacf071cc5a69faf28a63354b70578a3a9bcef29a928ac11c2468570bcac21d4d27af78a3bc1b00c25cda39b6`define QY0 381'h9385f2a6f2b6449ecc293f9fc4310e38b0745328b1732c619fbb8760801e13102ad3015aa92253d833cee0efa4cd993`define QY1 381'h1313ed4fe3934a5459c83660403bf785af03669baae7d60d5352b9b7bd78da012e52a668be24e635b04e4913b7cdf429`define QY_0 381'h10c8b2bfca5482505e5913bc47089bf3d9700652686ddff94d351a2aeeaf14f31bfecfe906c1dac236c211f105b2d118`define QY_1 381'h6ed249a55ec9c45f1537156030fb551b573e4e9489d3cb213de18e939381c22f0595995f32f19ca09b0b6ec4831b682`define TX0 381'h10b8501b92fe9329d24e30191ee6b5d10034a5eedfa61f71daaa1975e1b40b7c91a33c5021eff7f29fe39f429fa0a269`define TX1 381'h4ec8b6dacf071cc5a69faf28a63354b70578a3a9bcef29a928ac11c2468570bcac21d4d27af78a3bc1b00c25cda39b6`define TY0 381'h10c8b2bfca5482505e5913bc47089bf3d9700652686ddff94d351a2aeeaf14f31bfecfe906c1dac236c211f105b2d118`define TY1 381'h6ed249a55ec9c45f1537156030fb551b573e4e9489d3cb213de18e939381c22f0595995f32f19ca09b0b6ec4831b682`define TZ0 381'h5feee15c6801965b4e45849bcb453289b88b47b0c7aed4098cf2d5f094f09dbe15400014eac00004601000000005555`define TZ1 381'h0