`define PX 446'h19ca7f22d0bea5a5d368f623f0b1ae768dd06d03d82fdfda52fccb60bbe3aa1b276d14bbef02169fbb3208b84d83830516fd0d0b75916f43
`define PX_ 446'h231461d858073f8f4ca6cd2574f927c972c537b3b1d31e57bc78daeafee36be75ae15907f338b74e9bbc3c7077f032c71a1ef31b351f3b68
`define PX3 446'h10809c6d49760bbc5a2b1f226c6a3523a8dba253fe8ca15ce980bbd678e3e84ef3f8d06feacb75f0daa7d5002316d34313db26fbb603a31e
`define PY 446'h184a0369a8f205b05d7501d110bd3f10f5e1eb013cc28e98bd6b5ca403f84542c566c9c07dab1aef1f39001221d8cc13d32c959037adf72e
`define PY_ 446'h2494dd917fd3df84c29ac17854ed972f0ab3b9b64d406f99520a49a7b6ced0bfbce7a403648fb2ff37b54516a39ae9b85def6a967302b37d
`define QX0 446'h28dc6efd79f87ad77f2d784840970f83d53dd00f9cef017123817c2dba543781a77cf694dc4d9025a4959a608e2145520d3589222b67c8c0`define QX1 446'h3ae58e4c4241175f60a731494ffe3a4901c7742683c82b075dbaf98fb74ef72428130a6949e93a19229456a8e72b309f2bc11720be4b5b03`define QY0 446'h347440d7f2c3ba0687cbd18ec8f8ed6e42afcb33973d629ac90ba67019d2ce8f130b49579dc101c2436b90706aa89751eb2f8065eed06afe`define QY1 446'hf2f313a9977ab11dfa853c4bcc40aa91f6ca76b34d31b5e6236057d628d6be8a55490cfb57950575ab4317502e517a54a872f7d0aa73546`define QY_0 446'h86aa02336022b2e9843f1ba9cb1e8d1bde5d983f2c59b974669ffdba0f447736f43246c4479cc2c1382b4b85acb1e7a45ec7fc0bbe03fad`define QY_1 446'h2dafafc08f4e3a2340676f84a8e6cb96e128fd4c552fe2d3ad3fa0ce5839aa19dcf9dcf42cc17d96fc3a13b3c28e9e26e694d0a9a0097565`define TX0 446'h28dc6efd79f87ad77f2d784840970f83d53dd00f9cef017123817c2dba543781a77cf694dc4d9025a4959a608e2145520d3589222b67c8c0`define TX1 446'h3ae58e4c4241175f60a731494ffe3a4901c7742683c82b075dbaf98fb74ef72428130a6949e93a19229456a8e72b309f2bc11720be4b5b03`define TY0 446'h86aa02336022b2e9843f1ba9cb1e8d1bde5d983f2c59b974669ffdba0f447736f43246c4479cc2c1382b4b85acb1e7a45ec7fc0bbe03fad`define TY1 446'h2dafafc08f4e3a2340676f84a8e6cb96e128fd4c552fe2d3ad3fa0ce5839aa19dcf9dcf42cc17d96fc3a13b3c28e9e26e694d0a9a0097565`define TZ0 446'h3211f04d73a1acadff03cb69a5529bfff6a5b4875fd01cdf08a59b44538e9fd7db1923c1dc53211a911bad73a8c4a33cee3ffd9554f5555`define TZ1 446'h0