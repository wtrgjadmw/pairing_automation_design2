`define PX 381'h15c0fc57dee16c62760e8ba236b44029a96f45fd751deaf8700e90b19b8c2cd34603ff8bf82ddffe7715b0f21faa2183
`define PX_ 381'h44015925a9e7a37d50d1c140c976cadbb0805877e6727c6f72241ef5b24c950d8a80072b926200142e94f0de0558928
`define PX3 381'hd40d13329a477f2cbf4537a1d8566ce335f3aee784f9b6a81ca0cd2e5429a3194b3fea685e19ffbf14312d65eff0f33
`define PY 381'h11b83311edf1046db0b4da59dfaf573ea9001a38423b35ea3c29af87050f7e9064afcc627df79fb1ab94f27aa19caef9
`define PY_ 381'h848ded84b8ee22c9a66cd5c639c5598bb77314cb149dcd52b072319f1a17793b9fc339c335c604e0e6a0d855e62fbb2
`define QX0 381'hb03232486a179aedecf6ec630c66cd73129333a34795dd34351276a7c55cb0167ebf64d0f692c35ebe51f440528142
`define QX1 381'h15b312b0d98c0ab230ab9b6a90bb724a6ebccf7d474c047c74dacdbbd555879bec5518b2bc98ac184034780eb3c43ec1

`define TX0 381'hb03232486a179aedecf6ec630c66cd73129333a34795dd34351276a7c55cb0167ebf64d0f692c35ebe51f440528142
`define TX1 381'h15b312b0d98c0ab230ab9b6a90bb724a6ebccf7d474c047c74dacdbbd555879bec5518b2bc98ac184034780eb3c43ec1

`define QY0 381'h690c42c5e30150333c15f1c4ef0cfea309bc99e6aa2eddbd6c90555d2ed89f452da9f43981bd38b380e215f0c091434
`define QY1 381'h4a59a9173abc051a6466000dcf10ef89bb814fa779856bf3dbbcfe16652bc3886eac4e11b8d0c3b8cf7ff925bec8b61

`define QY_0 381'h13704dbddb4fd197175a4899f45adced33db81e688e224e39067cd4b23c36c2fcbd160bb19382c7481f0dea0f3f69677
`define QY_1 381'h155b7758c5d42648a4d547b5665a9ddec8bf368a7becbc00297502bf905e39eb97c13b1d95c6f3c42d07006da4131f4a

`define TY0 381'h13704dbddb4fd197175a4899f45adced33db81e688e224e39067cd4b23c36c2fcbd160bb19382c7481f0dea0f3f69677
`define TY1 381'h155b7758c5d42648a4d547b5665a9ddec8bf368a7becbc00297502bf905e39eb97c13b1d95c6f3c42d07006da4131f4a

`define TZ0 381'h5feee15c6801965b4e45849bcb453289b88b47b0c7aed4098cf2d5f094f09dbe15400014eac00004601000000005555
`define TZ1 381'h0

