// for wrapper -------------------------------------------------------------------------------------------------

// modes for the wrapper
`define I_INPUTMODE_SIZE    2
`define REF_RESULT                       2'd0
`define INPUT_COORD_CORE                 2'd1
`define EXEC_CORE                        2'd2
`define INPUT_CMD_CORE                   2'd3

// modes for the calculation core -------------------------------------------------------------------------------------------------
`define MODE_SIZE 'd4

// `define MODE_PDBL_FIRST 4'b0000
`define MODE_PDBL 4'b0001
`define MODE_PADD 4'b0010
`define MODE_PMINUS 4'b0011
`define MODE_SQUARE 4'b0100
`define MODE_SPARSE_MUL 4'b0101
`define MODE_CONJ 4'b0110
`define MODE_MUL 4'b0111
`define MODE_FROB 4'b1000
`define MODE_INV 4'b1001
`define MODE_MUL_CONJ 4'b1010
`define MODE_SQR012345 4'b1011

// for command buffer -----------------------------------------------------------------------------
// modes for the core 
`define CMD_SIZE   `MODE_SIZE + `RAM_ADDR_SIZE * 3

`define CMD_INSTTYPE 'd1
`define inst_ML 'b0
`define inst_FE 'b1
// for RAM -----------------------------------------------------------------------------

`define RAM_DEPTH 114
`define RAM_ADDR_SIZE 7


`define RAM_PX	    `RAM_ADDR_SIZE'd0
`define RAM_PY_	    `RAM_ADDR_SIZE'd1
`define RAM_BT0	    `RAM_ADDR_SIZE'd2
`define RAM_BT1	    `RAM_ADDR_SIZE'd3
`define RAM_PX_	    `RAM_ADDR_SIZE'd4
`define RAM_PY      `RAM_ADDR_SIZE'd5
`define RAM_QX0	    `RAM_ADDR_SIZE'd6
`define RAM_QX1	    `RAM_ADDR_SIZE'd7
`define RAM_QY0	    `RAM_ADDR_SIZE'd8
`define RAM_QY1	    `RAM_ADDR_SIZE'd9
`define RAM_QY_0	`RAM_ADDR_SIZE'd10
`define RAM_QY_1	`RAM_ADDR_SIZE'd11
`define RAM_TX0	    `RAM_ADDR_SIZE'd12
`define RAM_TX1	    `RAM_ADDR_SIZE'd13
`define RAM_TY0	    `RAM_ADDR_SIZE'd14
`define RAM_TY1	    `RAM_ADDR_SIZE'd15
`define RAM_TZ0	    `RAM_ADDR_SIZE'd16
`define RAM_TZ1	    `RAM_ADDR_SIZE'd17

`define RAM_XI10	`RAM_ADDR_SIZE'd18
`define RAM_XI11	`RAM_ADDR_SIZE'd19
`define RAM_XI20	`RAM_ADDR_SIZE'd20
`define RAM_XI21	`RAM_ADDR_SIZE'd21
`define RAM_XI30	`RAM_ADDR_SIZE'd22
`define RAM_XI31	`RAM_ADDR_SIZE'd23
`define RAM_XI40	`RAM_ADDR_SIZE'd24
`define RAM_XI41	`RAM_ADDR_SIZE'd25
`define RAM_XI50	`RAM_ADDR_SIZE'd26
`define RAM_XI51	`RAM_ADDR_SIZE'd27
`define RAM_ZERO	`RAM_ADDR_SIZE'd28
`define RAM_ONE	    `RAM_ADDR_SIZE'd29

`define RAM_A	`RAM_ADDR_SIZE'd30
`define RAM_B	`RAM_ADDR_SIZE'd42
`define RAM_C	`RAM_ADDR_SIZE'd54
`define RAM_D	`RAM_ADDR_SIZE'd66
`define RAM_E	`RAM_ADDR_SIZE'd78
`define RAM_F	`RAM_ADDR_SIZE'd90
`define RAM_G	`RAM_ADDR_SIZE'd102

// constants -------------------------------------------------------------------------------------------------
`define WORD_SIZE 'd1150
`define CHAR 1150'h39ef8b0000000000000bf301780000000000183380205001ee62800407b7a7590054f8ee04232eb06ee5aaa303908a651e230b8edc30861ef21c6df205d4fc8255bb46374c2a4afaba7fcb4ad0a05e8b00d7f54e6f78648c4d049d98d9575a0a520cf194d8c992014bb5886e2441a655668679e770013982d008555f4d5556200018c00009aaaaaaaaaadaaaaaaaaaab
`define CHAR_INV 1150'h22710f988516275bf316da7732c9fef8b657c67acec198be551f886d9fa08820164b41c6908179b0d381950dfa32b7a43d2b74e48023103e93ff03b7e59f208322582a9b716170a20e31ccaf7c2c40ee48e1fca77fd3e16aac0aa02bb1f2cebf003c8d5c4965a82ebf8a0347373f17e77dcd914b00470f59441dff5f20002df000debfff640000000001affffffffffd
`define INVERSION_INITIAL_VALUE 1150'h165a0d4fc86cf463ff78aff2fa7f0955fcba6e9bab32009bdda1d36944a8f4522839e14a075ca7c320c0012ae5844942f5ac742aa818b5391cd58addc65999b37b4009cf39bce67f9f6ebae43e82d1a7b5214c3d286b013e4ee67c68a314e5478807d8e1ea08c5599b7bca110c485e13f65be8ea59fff57d555a1c1c9c7bd68ec4cd91ee825339bbe61cf27b2aded3eb
`define CHAR_3X 1152'hadcea100000000000023d904680000000000489a8060f005cb27800c1726f60b00feeaca0c698c114cb0ffe90ab19f2f5a6922ac9491925cd65549d6117ef5870131d2a5e47ee0f02f7f61e071e11ba10287dfeb4e692da4e70dd8ca8c060e1ef626d4be8a5cb603e320994a6cc4f30033936db65003ac887019001de8000260004a40001d0000000000900000000001

// parameters for twisted curve (Ep2)
`define BT0 1150'h2b506ffffffffffff7c8eefd7fffffffffef5c97e9c8feac1c47fd3ab1bcf2cfc594dc5d27cfe6b3c21aafed8ca0da7b47e80dc89ea3cab98c74699bfd9266650f3fb9fba2ec739fc8243c9091bf006f6b875a135d3adf8b0cd3a6ea93f218e79719e9aaf56b9f1bf332344712dda549838c30e2ff287610fa454e7ad554c9ffeefbfff95aaaaaaaaa89aaaaaaaaaa7
`define BT1 1150'h61074fffffffffffff40cfe87ffffffffffe7cc7fdfaffe119d7ffbf84858a6ffab0711fbdcd14f911a555cfc6f759ae1dcf47123cf79e10de3920dfa2b037daa44b9c8b3d5b505458034b52f5fa174ff280ab190879b73b2fb626726a8a5f5adf30e6b27366dfeb44a7791dbbe59aa997986188ffec67d2ff7aaa0b2aaa9dfffe73ffff65555555555255555555555
// // constants independent from elliptic curve
`define ZERO 1150'd0
`define ONE 1150'h61074fffffffffffff40cfe87ffffffffffe7cc7fdfaffe119d7ffbf84858a6ffab0711fbdcd14f911a555cfc6f759ae1dcf47123cf79e10de3920dfa2b037daa44b9c8b3d5b505458034b52f5fa174ff280ab190879b73b2fb626726a8a5f5adf30e6b27366dfeb44a7791dbbe59aa997986188ffec67d2ff7aaa0b2aaa9dfffe73ffff65555555555255555555555

// Frobenius pre-calculated coefficients
`define XI10 1150'h2799e9b07192faa26b628d10c5d6ef6907c540ee96f61b76cb91b933cd38873cfc77c233b1e4e8dc5ed6dd488fcf213350c081aac290d549ccdb1071d120013f32bff07606d4f7c4498f2ea04e54183955a01ba805e516dd5725fb84a8eb78718d6787c33d2d0e0752440a9611c62522333164c5929f40ea63b53416bca06959a1acaae3653d7c3787566a73a28b5252
`define XI11 1150'hf95d2ef0f52b182f222b4dca1d94ae2e056dbd959f0202149591a0f69d8d62acb342538ff7d79d180255b33f8fd6fef9cb4cf04a1479d76d691b9b07ded98c07b3b72520ee84ab2dad8dc273b542e87c16b14b5a08c0177eeb5d5a1d20d38e803f0f7dc089d0d77aeba4d2655d7f555923ddc9d8dceacd80eb69be9c4355f65d370705cb370436d9cccc9b3a86ba7e9
`define XI20 1150'h247901549a7ba9ef2eb7278b8ba1c02a1d95de75df925e62294cfbb243725c3dd92c96120f1b0b9a2256c5594aa5d4cf393deb9c63bb55495675788d3d5cbc7ac97b1839bde295a987ac92e844bc01d30099723c8e49b5304ac94ee8c4cdd9199045c838cd9e99eee5012aceeaccf20a5c132dee1c3dd43201fc0b40a020268ae9353e709ef98ddda672116eeda5ab28
`define XI21 1150'h2c653568ed23bb7bb59a52eba836e6ea87f391a764526eded632c83f3a8539079049f54bec049e458987bc4f966ec509744b6cbe1b0644d1ce36710d19536b4c499615eb4d0560bf8badd8a8b7451b2d9cd881f60e48d9596caeeb9c83b605c289dbccd3d163d894c80d6e5d9c8e107253bd68495abc156778b7b4ea9da890629a35d9debca816088bef9946004a6bf
`define XI30 1150'h93230635b4f31267eb1364af3dc2669c42b8f76476d0c7362655cc20475d5b18f1f40fdf49660d5af3731edbd39b1fdac413f652023d8afe19e0d35f3d6131fafe03335b12007c7bb1c389ed4d3de7cef140963d5e417655361c33eb6f6428a32ee1bd9ed2c2795825b248e1b2d40ea0d534d29804036f25115ec6277b566b824b43225590ddcea0c2142f388a39298
`define XI31 1150'h220658e19117eb80f2e02bec0e998021a9b3826b4a222c7fe9931f9024e2b19696e390fd89bc99a8694248a660b069839c696e646535f0bfde1016298087c2ba8906b9e19f1602d2949a6ae97fa6525655f06897eb708568f4cd02da4c473f5bab4024ee6aeff9d5cbd9e51eeb82e2cf1eba89b79280ebf45ad2e6795fc0ad116ef1357570dff679cea1c2d8abb90f45
`define XI40 1150'h35c1002805b395aff6343a7d654f22d1492d191977537c05ed13b3d214ef56fc4ddf5d084caf9160c99e35fd8ddc8924e0c656acb4099b9ba4fa37cf946727cb0870f8de6ebcb5b5d2cec82c677522821d6125bfbc12a455842ccb59f7e3567ab817acd5680ac1b10a33ea59e07b8e431706cb0753d38e2b5aed973cf30a0b53e270bec59de4f61b782c8147c1b4219f
`define XI41 1150'h184e1fac968a4f974d6c8989e432d69bacd83c1a67723210995960e4884612372e67bc6550b3d2f8b2f7d65a3fa42e5b03216891140a2883de065c77020f5fa36ca061f598de97f6cc816a6ee9df36621c53a2dc25ceea58917442f0c7308f60ced936aa7a0fd1fd5dc0d5f32aa7b9b7a5f0f9bda3add5bf4f8645fd7429207d8ec1f5ebc8880c9b3cdbe21f6bdc2659
`define XI50 1150'h188a075517256bfc120172a803f79cebf7210d087eb5f99ded42ced6579f0c14d23d60e8834c8a279dfd37c7cc6e6f666b96212433425d26b69c8dde119fd093525df51eec727d48cac0bce5954d8ede778ddb6462d7be7c9e47147a34c9f0b12920424ebde16be2ed09afc8253124ce963ec7fc9c72cd319cee83ea92701fc2c575d9817341e972d7c13b7d6487f102
`define XI51 1150'hf5654d952122494ad859653599e25e25934ab9311cdfc3361671aeff4fcb41156ab0861f020667aacfc3b4219b525eb7580994087505fa8cd7d29b0c551fb1e6d4a08b8afdd8d79b59433077be34c4f4891c91bff3eb329016024e399a15795547bd56962f3fa73579c2570a3465e83deed1dbdf370946dccadbc3f955c1426e282221f0b770144c65cf31518adea22
`define CMD_MEMDEPTH_ML 584
`define CMD_MEMSIZE_ML 10

`define CMD_MEMDEPTH_FE 1013
`define CMD_MEMSIZE_FE 10

`define CMD_MEMSIZE 10
