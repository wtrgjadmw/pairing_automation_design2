`define PX 638'h251ae6f1843461ce31a2e2b50873a82d13ea5d6f9a77f6ad541dc0e4c5761e086091830e03198baf6326107c09b366ed96d58d4d4d4903248a00b0244449b7e1dfc127f77866ff718816f1a59396e2a1
`define PX_ 638'h179d8173b8fba971b65d32a0455eb583e8177f6efb5c0952ac455ad87ca0f6f8d8c3d24752391050f94fc646a14c9912692a7d7a48b7cf8720a9fa866660f2b20b32d7089243ab392293b9052b141d6a
`define PX3 638'h32984c6f4f6d1a2aace892c9cb889ad63fbd3b703993e407fbf626f10e4b4517e85f33d4b3fa070dccfc5ab1721a34c8c4809d2051da36c1f35765c222327d11b44f78e65e8a53a9ed9a2a45fc19a7d8
`define PY 638'h17fd7428a41951eff2d9522252aaedb48004b06f468251723f870917b40f9fe0973eec40e759fc68da0de54ad1cfa7aeee1919104b090e9b02de07ac0eb7a964c2cb4ccff5fa731b43a117fe222f3757
`define PY_ 638'h24baf43c9916b94ff526c332fb276ffc7bfd2c6f4f51ae8dc0dc12a58e077520a21669146df89f978267f177d930585111e6f1b74af7c410a7cca2fe9bf3012f2828b23014b0378f670992ac9c7bc8b4
`define QX0 638'h3184f22cd47d936ad263912e72bf659c71f8121b966eb0dba79c2d6ecdd851e11951adf85ca47f74b94a8dae92815ebca44deacaf02d99ec8c305000f5539ab116d2909459d112fd5625b6530200733b`define QX1 638'h360fc1eeaacef2aa432bb313d302e6f71e5320b47747966f6b4b36266edded8d434f4b8067fc5f02a99bd087523f4ad3ae6400597a7b33739462e896831b0a4e7bf94cdf2240bcafac8c827b3f2707f3`define QY0 638'h394d090243271a3fd607f4631d8ef07bb58241d2d03a8c9ae801d9f76f223ba0e6429acaf4b4d314bb5edddd4b76201f9af5f6fea08111b0a32bf75b0affed0639c7a3697e56a13a62fadec05c356b06`define QY1 638'hc7d30113b28fc4758a4f59325b966c59c444eb1326a1d85087f5983f523cc8aa385765c3ffd3b6aa445757c50037fe499f71de126b5639df0ba17d5c11193c1a46b98bb87f55077379b8b5859821607`define QY_0 638'h36b5f62fa08f10011f820f230436d35467f9b0bc5997365186141c5d2f4d9605312ba8a609dc8eba116f8e55f89dfe0650a13c8f57fc0fb077eb34f9faabd8db12c5b968c54097047afcbea62759505`define QY_1 638'h303b385402070ef88f5b1fc22818f6eb5fbd8e2d6369e27af7e3c2394cf3487695cfdef915556095b83061465afc801b6608ece66f4b6f0db9f092d4e99916d24688664482b55a33730f1f526528ea04`define TX0 638'h3184f22cd47d936ad263912e72bf659c71f8121b966eb0dba79c2d6ecdd851e11951adf85ca47f74b94a8dae92815ebca44deacaf02d99ec8c305000f5539ab116d2909459d112fd5625b6530200733b`define TX1 638'h360fc1eeaacef2aa432bb313d302e6f71e5320b47747966f6b4b36266edded8d434f4b8067fc5f02a99bd087523f4ad3ae6400597a7b33739462e896831b0a4e7bf94cdf2240bcafac8c827b3f2707f3`define TY0 638'h36b5f62fa08f10011f820f230436d35467f9b0bc5997365186141c5d2f4d9605312ba8a609dc8eba116f8e55f89dfe0650a13c8f57fc0fb077eb34f9faabd8db12c5b968c54097047afcbea62759505`define TY1 638'h303b385402070ef88f5b1fc22818f6eb5fbd8e2d6369e27af7e3c2394cf3487695cfdef915556095b83061465afc801b6608ece66f4b6f0db9f092d4e99916d24688664482b55a33730f1f526528ea04`define TZ0 638'h347979ac2cff4c017ffeaaab22da24f03fe23216a2bffffff9ce442bde8eafec6aaaaaaaaad63ffa38a293d54fffffffffff53869ff2d54555555555555556c150c00fff5555555555555554154fff5`define TZ1 638'h0