`define PX 509'h125e89836ae1ebab233be267497f2091b03f2f85e215a02e6aa54fdbfb4a8f402225306a23aaef4c9909ccafe9878217f94923d42eb96dffdcb95ed0fef4d034
`define PX_ 509'h2f6cd7c9457def0d9b2104db041cc651b4b98c37b02de5dc844b127e4c6017b40495555586db1a436c18fb0883351baf51a99333fd42500c483b2bcb9cb0277
`define PY 509'h11f2299602e0a2db8233f55f0dd60ffd44a076f2edd36c9c063d89228a3e2b4bd4acfa0dff0ffd1f04a831bf784d6239699bbc63ef0f135d7fc66b8f07b22cb9
`define PY_ 509'h3632d69fc5927c07ab9fd55ebeadcf986ea51566f4511f02cac77e155d2656f8dc18bb17d08a3d1cb232aa0f96d719984c800a37f7e7fa32176a5feb10da5f2
`define QX00 509'h45734dbcdf2412672a2f6b31766747f92e99a09328c8f62ddbbac12e1d6e8b3f8c9ed26ba1b15a4dba1d5b6d43be666831879ce38d601c51bbaa096f016b1c7
`define QX01 509'h134d1f64cf5f707d4d4110945773ca8a8fcbe031708e8123b95c001596b08b3723d41541408665ebfd0463e6a2fe67f5cb782366940f1fae7cf184ccfa89b557
`define QX10 509'h1373b923cb62bc6595c92a9777219765f56f7bfda1cca7ad086c83a8099654e07f06f2cf6a40cd1d1b7a5fa6cd8e704cfa84926794f0bca79bf8cde6bf1e83e6
`define QX11 509'h194cb42691c401c0b3d635d4d2cf62a1481af2efca3c388cb0c2cbcec9970579ca6b75c7402e8a714f448a0873f3c200eae45b1cf4d8e4f1c54ebb0200dd27d
`define QY00 509'h3dfbf874af39807b76429fe5c4818e5a83e392583a9ec39b22a10b138774dc0f593b080537fd9fe9a539a298dbf77750d2dea03d43f076ce94e4f168ba56ab0
`define QY01 509'h117176e910de242d2d3be0c9edc218292d3e0037e32ec43efc46858cfafcf4429eae50f90fa4572487c532a59d785f54180849f3cf9dca3632e190c9f9cff443
`define QY10 509'hacbe80c5817a708aca98a1a9983e7ec2cef0e602e09b6cd4a362fb009665a04bfc2357d1fa02225261857595fe395a76e15f606846576da440bb9dc7e582c53
`define QY11 509'h7f8ee90e7816b48cd858ca0a8dcae1f0ac5b3ef37274fb665c95c65b4d2f2d85fa3660dd2b521beab0d15b2a40656c16eeec147bcc6acedbabc5c95ed59e5ae
`define QY_00 509'h11759778b44632944589c8b69d78d411234c8f23d96e925280bff052a79942fa6cdad53f2898c6f23577c236e3fb5c5de135d3039a4e8b93b7eec2772d1a67fb
`define QY_01 509'h3e3e016ee5ba66ecfb211eb0bfed4cd9e4cc81179e9ba4d36a37b76e5139c78c3c034c66c7449cc480629bad442747ed65b73139eefc8ca6e5b80c3beefde68
`define QY_10 509'ha896ef3a72223935044689a603d050a9e9bb9e92f0ec7bee8b3d153d6aa36b6a2ac50425c787ecba9b3050711d73e2b804dc700ea281c265d3157b13a67a658
`define QY_11 509'hd5c686f17b85f532f68661450e43ed7c0c5145a25f12ed5cd20a49e2b3d9de302cb1fb1a9637f3224be46adcdb47d117f74fbbfb1c6e612e680b4f7cb65ecfd
`define TX00 509'h45734dbcdf2412672a2f6b31766747f92e99a09328c8f62ddbbac12e1d6e8b3f8c9ed26ba1b15a4dba1d5b6d43be666831879ce38d601c51bbaa096f016b1c7
`define TX01 509'h134d1f64cf5f707d4d4110945773ca8a8fcbe031708e8123b95c001596b08b3723d41541408665ebfd0463e6a2fe67f5cb782366940f1fae7cf184ccfa89b557
`define TX10 509'h1373b923cb62bc6595c92a9777219765f56f7bfda1cca7ad086c83a8099654e07f06f2cf6a40cd1d1b7a5fa6cd8e704cfa84926794f0bca79bf8cde6bf1e83e6
`define TX11 509'h194cb42691c401c0b3d635d4d2cf62a1481af2efca3c388cb0c2cbcec9970579ca6b75c7402e8a714f448a0873f3c200eae45b1cf4d8e4f1c54ebb0200dd27d
`define TY00 509'h11759778b44632944589c8b69d78d411234c8f23d96e925280bff052a79942fa6cdad53f2898c6f23577c236e3fb5c5de135d3039a4e8b93b7eec2772d1a67fb
`define TY01 509'h3e3e016ee5ba66ecfb211eb0bfed4cd9e4cc81179e9ba4d36a37b76e5139c78c3c034c66c7449cc480629bad442747ed65b73139eefc8ca6e5b80c3beefde68
`define TY10 509'ha896ef3a72223935044689a603d050a9e9bb9e92f0ec7bee8b3d153d6aa36b6a2ac50425c787ecba9b3050711d73e2b804dc700ea281c265d3157b13a67a658
`define TY11 509'hd5c686f17b85f532f68661450e43ed7c0c5145a25f12ed5cd20a49e2b3d9de302cb1fb1a9637f3224be46adcdb47d117f74fbbfb1c6e612e680b4f7cb65ecfd
`define TZ00 509'haaaa90000c6356403120d4b063f1309347537b6a2e78173cd15fefc1fef6f449d917a4083e75f0f3034a39f8e452c2d119c42f891726cff5ec2ee7247402d55
`define TZ01 509'h0
`define TZ10 509'h0
`define TZ11 509'h0
