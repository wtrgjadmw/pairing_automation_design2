`define PX 1150'heba940b8314fe6ff2a8025a0a632453afaee2776fc9b80a05f73295be7bae0c96e28a2878e3b5aa49cf4dd27dcd3a6d65e68d9a1631fca35096e3e358401ab5e02c9c907d98250bd57d632f2dd0d594112e18d3ea62a12591ffcc186605f1efb5e4c8557dd9cc497382e16edd1b754d63df7b8a2b139c224fb61e5d57feab8ea748a909d7f9b41b439e21724a2367df
`define PX_ 1150'h2b34f6f47ceb01900d63f0a76d9cdbac505135bc105697f7e86b4d6e493bf94c69726ec58b3f790625165cd085c34ff7b83c7df4c5fe897ba1858a0ead94e1cc758ea9a6ce9225eee502681ba2cf88f6efa9dc7a8515c366bb04d1807351681a9c28293f5aefc5b7d832a6ff4726310802a6fe5d44ed9d6080523701f556aa9158d016f631b0f68f670cb938608742cc
`define PX3 1150'h2c2fbc22893efb4fd7f8070e1f296cfb0f0ca7664f5d281e11e597c13b730a25c4a79e796aab20fedd6de9777967af4831b3a8ce4295f5e9f1c4abaa08c05021a085d5b178c86f238078298d897280bc338a4a7bbf27e370b5ff64493211d5cf21ae5900798d64dc5a88a44c97525fe82b9e729e813ad466ef225b1807fc02abf5d9fb1d87ed1c51cada6456de6a379d
`define PY 1150'h388b49db3fc982dc213e65f6d530a82364e1039327dfa04eae3ada84e6c44790645327db8916689a6918b92321105022e6e21803c5a8ae98f4a1ee6a7912936b379268852024167a80f4bb611c8fec9bd0636eacc24fde3e6aee57e08c804b47659afd97a9b28cc8b7ce3dc4fd77d93f53de963147e4057014e9deaad0d4fedb2326ca943e44fe531845599e33d633e4
`define PY_ 1150'h1644124c0367d23decd8d0aa2cf57dc9b1f14a05840afb34027a57f20f35fc89c01d1127b0cc61605ccf17fe2803a423740f38b1687d785fd7a7f878cc269171e28ddb22c063480398b0fe9b41071ef307486a1ad28864de21645b84cd70ec2ec71f3fd2f17053893e74aa926c9cd1612a7e3b6281d3412bb1e76b47c805744dcf1f56bcb65ac579265810c76d476c7
`define QX0 1150'h16258d52f49106c4b53771c2edf54e74d996499fc9c3f08a9f8a67fcc611b85ec3dcc9fb1c2daef8bb506f0716312f277e3cd38b34519147045d9ad9497b5a510a5590e6168fa29cca60ab9d0a87c40686b0750b7a1b9ea7319adb716a47d12c0bf314ff84cc64a5d7ad7479aa8212fdbf022e6b2688e92403771cd67d247c83c69846815fe26c755eba5a1d39c1b78f`define QX1 1150'h1552cc5f5fa7f75f8a89949b64765df9eb7e63fb3b4a4b9be52f442a22ba27364497c4a1419348b0fb423170d50b6c56bbea19b3c93a645d22236134e7ee5fd599cb65f1498d97d4ddba75e560b0291ccac7451b9aaa2dc0f0610ae64150268f85f5d4be5882508a2f5e10cc3ac1cb2398bcf4878a946eae14682a582a5fb58c1982589a900e6308f72d7eed6ecde635`define QY0 1150'h118f8d42b9ad17da54bef323852fcd68e3e8c700576414cfae7167c08ad3d1af081d8ca60764aed98fea9b231011166ecebb8e564968ebc519d9465346784873a327874b6a3fd49dee82a924fed7088d4834a095f8aca8e82235c5fd263405fc6040dde3818f2e8cb01214051105401a44e15f740673162ddc2b79ebcbb0d98ff207199ee5056c606f9457973c6b6da9`define QY1 1150'h97f285210c4fdf63ecf133f35924948388614fc88ff65ee8aac8a5990420c378e4d1d089a26d0f17e7ce8e5d663319e8a111e180a880e51823155b62d1deec5547205a3fad6dda8f548a11b61484ad5dd3c6a74119e474c3102570fea5e15ce2a0ee5c64ded526fa3b5dea29cbc144d6d3a6ed1b066340159341ddd79297d003eb99ab980c614339e5c5def695e1877`define QY_0 1150'h285ffdbd4652e825ab4cffddf2d032971c17513328bc3b323ff118437ce3d5a9f8376c47fcbe7fd6defb0f7ff37f73f64f677d3892c79a59d843279ebf5cb40eb293beebe1ea765ccbfd2225d1c955fdb8a354b876cbbba42aced79bb323540df1cc13b1573a63749ba37469133c663b21a51a73698e2354f3dcdb7381a47c900e11a66124a53e4a3b1683136e3f3d02`define QY_1 1150'h307062adef3b0209c13cdfc2426db6b7c77a0336f720ea1363b5f5aa77759b217207dbe569fc5dbef068c1bd2d2d58c69411ed76d1a877cd6feb183bd8b70dbd0149409351536d51c5372a2f6f5813b5239b8ada5dda1d401c024688eef9443c27fe0bce8adc3f91a7ffa9cb87859207f94c0b15bf9b058176d43781d42bd91fc15f254688e496770c4e7cbb414c9234`define TX0 1150'h16258d52f49106c4b53771c2edf54e74d996499fc9c3f08a9f8a67fcc611b85ec3dcc9fb1c2daef8bb506f0716312f277e3cd38b34519147045d9ad9497b5a510a5590e6168fa29cca60ab9d0a87c40686b0750b7a1b9ea7319adb716a47d12c0bf314ff84cc64a5d7ad7479aa8212fdbf022e6b2688e92403771cd67d247c83c69846815fe26c755eba5a1d39c1b78f`define TX1 1150'h1552cc5f5fa7f75f8a89949b64765df9eb7e63fb3b4a4b9be52f442a22ba27364497c4a1419348b0fb423170d50b6c56bbea19b3c93a645d22236134e7ee5fd599cb65f1498d97d4ddba75e560b0291ccac7451b9aaa2dc0f0610ae64150268f85f5d4be5882508a2f5e10cc3ac1cb2398bcf4878a946eae14682a582a5fb58c1982589a900e6308f72d7eed6ecde635`define TY0 1150'h285ffdbd4652e825ab4cffddf2d032971c17513328bc3b323ff118437ce3d5a9f8376c47fcbe7fd6defb0f7ff37f73f64f677d3892c79a59d843279ebf5cb40eb293beebe1ea765ccbfd2225d1c955fdb8a354b876cbbba42aced79bb323540df1cc13b1573a63749ba37469133c663b21a51a73698e2354f3dcdb7381a47c900e11a66124a53e4a3b1683136e3f3d02`define TY1 1150'h307062adef3b0209c13cdfc2426db6b7c77a0336f720ea1363b5f5aa77759b217207dbe569fc5dbef068c1bd2d2d58c69411ed76d1a877cd6feb183bd8b70dbd0149409351536d51c5372a2f6f5813b5239b8ada5dda1d401c024688eef9443c27fe0bce8adc3f91a7ffa9cb87859207f94c0b15bf9b058176d43781d42bd91fc15f254688e496770c4e7cbb414c9234`define TZ0 1150'h61074fffffffffffff40cfe87ffffffffffe7cc7fdfaffe119d7ffbf84858a6ffab0711fbdcd14f911a555cfc6f759ae1dcf47123cf79e10de3920dfa2b037daa44b9c8b3d5b505458034b52f5fa174ff280ab190879b73b2fb626726a8a5f5adf30e6b27366dfeb44a7791dbbe59aa997986188ffec67d2ff7aaa0b2aaa9dfffe73ffff65555555555255555555555`define TZ1 1150'h0