`define PX 638'h15f991ebd2849c8902483b04a33126eec7cee03a2845a308b2cf58fb2d39cde922ff87a82b5a792d32424b51eef701dd438e3a6c199edbcbcb72b90f093c70533bbff2ab6cee82530654e227f62f2664
`define PX_ 638'h26bed6796aab6eb6e5b7da50aaa136c23432fca46d8e5cf74d93c2c214dd47181655cdad29f822d32a338b70bc08fe22bc71d05b7c61f6dfdf37f19ba16e3a40af340c549dbc2857a455c882c87bd9a7
`define PX3 638'h5344d5e3a5dca5b1ed89bb89bc1171b5b6ac3cfe2fce91a180aef34459654ba2fa941a32cbccf873a510b3321e50597caaaa47cb6dbc0b7b7ad8082710aa665c84bd9023c20dc4e6853fbcd23e27321
`define PY 638'h15145fb2acc8b40893ff9b3c8d2962695f65d158afe75bbcf7fecc68c73704515a410e822a7c3b5507d866e577c70d5c4d2436aa6aa6057fec64a13c96942f570f3b0683f2f2a3568414f52b79ba438e
`define PY_ 638'h27a408b29067573754007a18c0a8fb479c9c0b85e5eca44308644f547ae010afdf1446d32ad660ab549d6fdd3338f2a3b2dbd41d2b5acd2bbe46096e14167b3cdbb8f87c17b807542695b57f44f0bc7d
`define QX0 638'h5fe3d09e2be654fd862a4ce349d4e76b602a66ec014fb46f1413a08d12607bbd64f59e835f22d7f2e7036c93c9f072a9123fcdc1311591b22fc2cc4eadc44387be9c1b614707d7716c6e1c3d685039a`define QX1 638'h3640a263cbd212429267aeeab006073ccbf9ae502c69bef907b3c2a86d333a8c181a39acde2c8ac1a6e9d8c3bf9c99157a3e64a0d33e849f8f7e0e8f18961ef626af425439399d4ee525c593830471c5`define QY0 638'h368264406ce32c7932998f2033de2cf4d5010408e0f3330d005cefe6cddf146bf75673f1ad0df060af853d417ff4310754d9e9a6435bfa02ca4b0ce5205e2bc363997ac2ebe33ed36e880738af9df950`define QY1 638'h1f7147bfef5b8a9d4c345bcd5e94258201ac8012f38a49de69389a3877f9111e47c0722e83781b933d1a8efebd189ce5c996c0e3532957433dc9ea917c29894217a83d9a3293dc09d8aa8085071d6bfc`define QY_0 638'h6360424d04cdec6b566863519f430bc2700d8d5b4e0ccf300062bd67438009541fee163a844ab9facf099812b0bcef8ab26212152a4d8a8e05f9dc58a4c7ed0875a843d1ec76bd73c22a3720f0d06bb`define QY_1 638'h1d4720a54dd480a29bcbb987ef3e382efa555ccba249b621972a8184ca1e03e2f194e326d1da806d1f5b47c3ede7631a366949e442d77b686ce0c0192e812151d34bc165d816cea0d2002a25b78d940f`define TX0 638'h5fe3d09e2be654fd862a4ce349d4e76b602a66ec014fb46f1413a08d12607bbd64f59e835f22d7f2e7036c93c9f072a9123fcdc1311591b22fc2cc4eadc44387be9c1b614707d7716c6e1c3d685039a`define TX1 638'h3640a263cbd212429267aeeab006073ccbf9ae502c69bef907b3c2a86d333a8c181a39acde2c8ac1a6e9d8c3bf9c99157a3e64a0d33e849f8f7e0e8f18961ef626af425439399d4ee525c593830471c5`define TY0 638'h6360424d04cdec6b566863519f430bc2700d8d5b4e0ccf300062bd67438009541fee163a844ab9facf099812b0bcef8ab26212152a4d8a8e05f9dc58a4c7ed0875a843d1ec76bd73c22a3720f0d06bb`define TY1 638'h1d4720a54dd480a29bcbb987ef3e382efa555ccba249b621972a8184ca1e03e2f194e326d1da806d1f5b47c3ede7631a366949e442d77b686ce0c0192e812151d34bc165d816cea0d2002a25b78d940f`define TZ0 638'h347979ac2cff4c017ffeaaab22da24f03fe23216a2bffffff9ce442bde8eafec6aaaaaaaaad63ffa38a293d54fffffffffff53869ff2d54555555555555556c150c00fff5555555555555554154fff5`define TZ1 638'h0