`define PX 509'h13681aafdfb5d016a0e1528e066854c7c91f092b681ac0e65c1a32310e96a278d8aae0c2fcb9c793956c1e6d0e32db963bee0c7d7291d1e2e056c72c506b16e3
`define PX_ 509'h1ed3c501f83fa855c0ca026f358982f026bbf1df4fdbda5d6cfced2d179ee4289c3a4fc7f5ed95d3a5f3df36387f83cb275b089fbfbc11dc0e64a616854bbc8
`define PY 509'h2021d1b0c8dace0ef7fee87f1770b3bd8ba0f7a11231251563521fdfc90e30d5fa5db731a640711db2b5d3c4780af3b40f57c20caf52a12606ebebb931fc7af
`define PY_ 509'h135339e4f2ac1dbb0d6e042d0849e1baf2d0b8cf4bf56c3adcb4df05e37fadae02c8aa4c61b499def49fff242a3a2497ad6e40e6a39868ee40ce52d225a00afc
`define QX00 509'hdd84c16d9d0722bbf84807fd17b26ed90bdad0353c10a16b4f2a92a492be904302381e813520c6ee43bd80dfbffee94cea163b11aad6014d6d2f7079bce4174
`define QX01 509'h9604ed78aba133ab55bfa4431d05ba2178d7ede856f36fa2bc6be6e5edfc9b8da02414178f07ced5ffd71f45a25ecb57b6c91363e4aaab6de006d06f46c91e5
`define QX10 509'h780b33e9b84a6aaf1a36a8cb3bf62abaf6c537feb489a9e0bfa17c7205f2e09ac884e8725a3056474ef1c4a96bc2a65fd832f4ce113f1d88fc73b4939e4d436
`define QX11 509'h96d393d966e3317c057fab977a238a7aa73281d2a23ee7b545bb470429decfab1da749df745e6a96b81118db3edda7a2e1b4986c96f25f2c7b4b0bb06af5849
`define QY00 509'h141996bd5d57b02684e82b2e0cb44b4148eab08353f5e005ecd9f85307087defc80785f9f3fda33d37358dfa96f6a09c3d3067c1917c4696327c24f05f840587
`define QY01 509'h3d48c1514c15fe80648634897da1c412b73ca65716f288a7af85ffb97a114dc47f226f38f89f36900e6327da18aeb44f08ebc771334ae14bdc77695e87804fc
`define QY10 509'h926fa3dc689761ad21b30195bad80702238f876777636239cc5e56b33b64a7559e54a87421652e4e558345d34af3d8e21f1e291def5a7a938fd43d72d614d38
`define QY11 509'h4ecadcdb69e4d8e022085859258b13ff18515b53599efdf7266da3bc7252af523df2ce8f94477548366c3a3ca144db007e479afa26def7c71ab16f6ddccc77
`define QY_00 509'h13bc042a1e21a757805c786ed0ca1b582a017c609229e86461008b0d90812cb9a66ffc5881afdb39895ce65dac43336b1335545dd114c6a6ec0ec9d593bcd24
`define QY_01 509'h1180caeaea786ab3f6a58f6c61e6d0b5a016fde3eba95601b7f1a108486f7bdf1a7c5ecbec8ead87cee529e2d02fe88dfdd500905b58e4ebe3759af7d047cdaf
`define QY_10 509'hc2e5cc238b054812ad2c29b9e136c86a951cfd2e5a2486896241b98ac5a464608893b383a024e0bea7328033d0b9644cc71da758f97eb57683fcdb68b5e8573
`define QY_11 509'h15068c2323cfe5c31ccbea5ca09b61e2cc7276ee09bedf8e3bc39360239e3e0c103092f0ec84597b8794f02635198ef7ede5756c7466b408da22601e4ae30634
`define TX00 509'hdd84c16d9d0722bbf84807fd17b26ed90bdad0353c10a16b4f2a92a492be904302381e813520c6ee43bd80dfbffee94cea163b11aad6014d6d2f7079bce4174
`define TX01 509'h9604ed78aba133ab55bfa4431d05ba2178d7ede856f36fa2bc6be6e5edfc9b8da02414178f07ced5ffd71f45a25ecb57b6c91363e4aaab6de006d06f46c91e5
`define TX10 509'h780b33e9b84a6aaf1a36a8cb3bf62abaf6c537feb489a9e0bfa17c7205f2e09ac884e8725a3056474ef1c4a96bc2a65fd832f4ce113f1d88fc73b4939e4d436
`define TX11 509'h96d393d966e3317c057fab977a238a7aa73281d2a23ee7b545bb470429decfab1da749df745e6a96b81118db3edda7a2e1b4986c96f25f2c7b4b0bb06af5849
`define TY00 509'h13bc042a1e21a757805c786ed0ca1b582a017c609229e86461008b0d90812cb9a66ffc5881afdb39895ce65dac43336b1335545dd114c6a6ec0ec9d593bcd24
`define TY01 509'h1180caeaea786ab3f6a58f6c61e6d0b5a016fde3eba95601b7f1a108486f7bdf1a7c5ecbec8ead87cee529e2d02fe88dfdd500905b58e4ebe3759af7d047cdaf
`define TY10 509'hc2e5cc238b054812ad2c29b9e136c86a951cfd2e5a2486896241b98ac5a464608893b383a024e0bea7328033d0b9644cc71da758f97eb57683fcdb68b5e8573
`define TY11 509'h15068c2323cfe5c31ccbea5ca09b61e2cc7276ee09bedf8e3bc39360239e3e0c103092f0ec84597b8794f02635198ef7ede5756c7466b408da22601e4ae30634
`define TZ00 509'haaaa90000c6356403120d4b063f1309347537b6a2e78173cd15fefc1fef6f449d917a4083e75f0f3034a39f8e452c2d119c42f891726cff5ec2ee7247402d55
`define TZ01 509'h0
`define TZ10 509'h0
`define TZ11 509'h0
