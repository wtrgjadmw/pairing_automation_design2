`define PX 315'h272409190897cadb98aba1af04e7b76677f15dd00e2566c48940c1edccdd6fb0410d2228288d8ee
`define PX_ 315'h24ff97124fd59a31a6c8f70f92de3397742ba3da197c473f98ad9bb75f00e076bd730dcbda72713
`define PY 315'h30d4b75165933e99143bc79055dc2bfc4cf85c0264f50cae8ee6d3b305e8369735f2b3cd82dc386
`define PY_ 315'h1b4ee8d9f2da26742b38d12e41e9bf019f24a5a7c2aca155930789f225f6198fc88d7c268023c7b
`define QX00 315'h17191cc8c571bd7dfacd0d47e0b22debae7cf1f30802cebc61d95aa4ac11fbc5e928b7b90ffcb96
`define QX01 315'h2b3179592438f93ba606f8f57e2101c53c1aa5252c8d709b0854c5e364390e1426738cf852aa221
`define QX10 315'h1834b8050ba6b271e23abc109d398998a1ad9837ccfe1e9a9dc8d67a9bbc7676d32ef6218aa5134
`define QX11 315'h1dd66aee1da974c6e5aef5be45ac5f00e75f1a3dd9d3e33307bc9726fc462f3cbb99d9364575cd
`define QY00 315'h15b0673b73e18e5fc7c2e4ea8c51f1977cb50c53acc080b176252a674e6b1a9353c3971ef869a53
`define QY01 315'h29ff47c749dd82f3128853b4a42cb87087f9772b7dc2a4abbd99a76877a0e04e90c9694162d24e
`define QY10 315'hb816dcc7cbe128d8fcb2bd4f59ad2ace4fc7a4e588c76a2e8b2058f7a12e123d4785c925a53504
`define QY11 315'h2dbd022ba26515a31322f2f29a1d1f912ae4a9ce9d71a7a5489a50f0c62b856e26daa8317eb60a5
`define QY_00 315'h367338efe48bd6ad77b1b3d40b73f9666f67f5567ae12d52abc9333ddd733593aabc98d50a965ae
`define QY_01 315'h4983abaee3cf8cde0e4c13834d831f76e39d6a376fc583b96614c32ea46442221573995fecd2db3
`define QY_10 315'h40a2325edbaf527fafa96ce9a22b18510720875bcf153761393c5815b1cb6f032a07d361a8acafd
`define QY_11 315'h1e669dffb6084f6a2c51a5cbfda8cb6cc13857db8a30065ed9540cb465b2cab8d7a587c28449f5c
`define TX00 315'h17191cc8c571bd7dfacd0d47e0b22debae7cf1f30802cebc61d95aa4ac11fbc5e928b7b90ffcb96
`define TX01 315'h2b3179592438f93ba606f8f57e2101c53c1aa5252c8d709b0854c5e364390e1426738cf852aa221
`define TX10 315'h1834b8050ba6b271e23abc109d398998a1ad9837ccfe1e9a9dc8d67a9bbc7676d32ef6218aa5134
`define TX11 315'h1dd66aee1da974c6e5aef5be45ac5f00e75f1a3dd9d3e33307bc9726fc462f3cbb99d9364575cd
`define TY00 315'h367338efe48bd6ad77b1b3d40b73f9666f67f5567ae12d52abc9333ddd733593aabc98d50a965ae
`define TY01 315'h4983abaee3cf8cde0e4c13834d831f76e39d6a376fc583b96614c32ea46442221573995fecd2db3
`define TY10 315'h40a2325edbaf527fafa96ce9a22b18510720875bcf153761393c5815b1cb6f032a07d361a8acafd
`define TY11 315'h1e669dffb6084f6a2c51a5cbfda8cb6cc13857db8a30065ed9540cb465b2cab8d7a587c28449f5c
`define TZ00 315'h33dc5fd4a7929af2c08b6741683a150213e2fe55d85e51fbde11a25ad421afd9017fd00bfcfffff
`define TZ01 315'h0
`define TZ10 315'h0
`define TZ11 315'h0
