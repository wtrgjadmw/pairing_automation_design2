`define PX 318'hca3ff498a4ad0337b6ed002e3cfd3947281a3713efff98d80821fbcddc7d43cdadaace655ffeffa
`define PX_ 318'h201ce66fa6c2cb399f5913423f15fdf47e44852d972121369c3d97dffe730b82257a49195a556ab1
`define PY 318'h16a93b3e69746de68ac9170acffac8c3ac412bc475c85cdece375c61773145255e86513d74918754
`define PY_ 318'h1617aa7ac7992d868ffecc3a52eb08c54484fcda6058bde54e885b3b65099a99a1cea4c23bc3d357
`define QX00 318'h8ea112b6dc3f7867056eaec3d712cecc850521e04117fcbd7a92123bdc8a3b7f03b989669a0a209
`define QX01 318'h171e096b4ad82b2772b4cb71faf6b81536f915a16e439ea83fd31a79b0de981fea1ed64e767ecdab
`define QX10 318'h51b033f6b56c3bdcbfc54fca0e962419f8aab8cf9dcdbe798107a0bc26375a29e333763875d283
`define QX11 318'h22bb87d3b7ff13b0220ffe3621d8c589a54390681e088e694a011d4a181ed6116d19b5c62451f455
`define QY00 318'h11eeeb84e29409026137dc82cfb57c2b53a19ef42c02144ba62d1bf13bdc08ea2223265219e627b9
`define QY01 318'h2b6d7eaaec6752997bc643aa7e61e598375165d888816fe78799d10d616566f54175268059f39d5a
`define QY10 318'h132aa9a9cc1e629c9a572b29430669b9bef664e821b61001076e6da887a6711dd6a8c3677ba85294
`define QY11 318'h25784ab870356e80a00e3655fd5208e73e6ce1e97d437273317ed4404717a2f09e30c0b558e20c69
`define QY_00 318'h1ad1fa344e79926ab99006c25330555d9d2489aaaa1f067876929baba05ed6d4de31cfad966f32f2
`define QY_01 318'h153670e44a648d39f019f9aa483ebf0b974c2c64d9faadc9525e68f7ad578c9bedfcf7f5661bd51
`define QY_10 318'h19963c0f64ef38d08070b81bdfdf67cf31cfc3b6b46b0ac3155149f454946ea129ac329834ad0817
`define QY_11 318'h7489b00c0d82cec7ab9acef2593c8a1b25946b558dda850eb40e35c95233cce6224354a57734e42
`define TX00 318'h8ea112b6dc3f7867056eaec3d712cecc850521e04117fcbd7a92123bdc8a3b7f03b989669a0a209
`define TX01 318'h171e096b4ad82b2772b4cb71faf6b81536f915a16e439ea83fd31a79b0de981fea1ed64e767ecdab
`define TX10 318'h51b033f6b56c3bdcbfc54fca0e962419f8aab8cf9dcdbe798107a0bc26375a29e333763875d283
`define TX11 318'h22bb87d3b7ff13b0220ffe3621d8c589a54390681e088e694a011d4a181ed6116d19b5c62451f455
`define TY00 318'h1ad1fa344e79926ab99006c25330555d9d2489aaaa1f067876929baba05ed6d4de31cfad966f32f2
`define TY01 318'h153670e44a648d39f019f9aa483ebf0b974c2c64d9faadc9525e68f7ad578c9bedfcf7f5661bd51
`define TY10 318'h19963c0f64ef38d08070b81bdfdf67cf31cfc3b6b46b0ac3155149f454946ea129ac329834ad0817
`define TY11 318'h7489b00c0d82cec7ab9acef2593c8a1b25946b558dda850eb40e35c95233cce6224354a57734e42
`define TZ00 318'h133f1a46cef26492e5381cbadd1a2e770f39d76129dee53be340486323c52040ffab0a004faaa555
`define TZ01 318'h0
`define TZ10 318'h0
`define TZ11 318'h0
