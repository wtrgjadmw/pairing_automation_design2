`define PX 1032'h5f766b8a8e6a296ce86b73483598427c51cc2026c4d47d5493e5f86078e7207b89eb5cc26dce475fea1193e55a001215fc6f54bb47cf85dc3e9a78495b5964bfea66c727ed3a57b2428c1828949940ad12b57a4ddf31522d0017a4719e31c2af9901c18d8dd9c626fb0229d3a61332eb884bc03cc5b05c53f27016391d6d11d839
`define PX_ 1032'h673835ca003c58e7c8a793167ccd1da75e00b8cc44ce1865bc20fe52a27ad8fae288f3f36a2f15505f546e4299a37252f6e0633669d156e9627b528af6ba85a3901e66c373379e244dd6fc56361e3bca22aadf073f2278d2876860f3c2ce3fb066e0e8fd1ccb8f4f5a532b7b0495cd14cd09bfc30a4fa3ac12e540718d3d98d272
`define PY 1032'h476cd84cb89257a3940fecc796c350ee88c5944f34a477df75985ea0e3951fbbc6e3cb4384d188cae2360db724c2ad892e4a23991cd2dd487382001dc16f235fd19ef5ab51233ff3984afd3c771873075b20db0b3fe7de6860a4cdee93116654f5b6bb6927b5d8700cb917483289f171da663f2e590b834505e6d8ab1efaadf75b
`define PY_ 1032'h7f41c907d6142ab11d0319971ba20f35270744a3d4fe1ddada6e981237ccd9baa5908572532bd3e5672ff470cee0d6dfc505945894cdff7d2d93cab690a4c703a8e638400f4eb5e2f8181742539f096fda3f7e49de6bec9726db3776cdee9c0b0a2bef2182ef7d06489c3e06781f0e8e7aef40d176f47cbaff6e7dff8baffcb350
`define QX00 1032'ha6956d27f52dc6f7460a7a97a5741f3b78d967e63f77a0b2e804e865e272cade37483ff1ccbf7092ded3f182434c3a528b123df309324a222d3df4d15f5fd0391d3f3a9b0458ebbabb62f0527fc93993d3cfa22c4ccb05e6a251512a9762a9b43ff301ba725bbb59639af50bd30865d6379700bbe99021736997d97deaa61a0288
`define QX01 1032'ha1e60a0f4df7a90eb30f2dc816893131194d296b2eb3c5479027ee25924d3dcb6ab2eb0bc380f1d7cf27c460b8eee6d62726c4b11344ba399fc7ff1ad487f5bbb7e632e2d44c019f69b8c692559c8cb28f4163c3119661f37b0cb22b13af8ada73cfc6fa132e20801dcb8ef907db5ed9a3f8b4312fb87070efb9461b84aa285bb2
`define QX10 1032'h1f842bd54a96d9a42b1d576b636d4ced5a61305ac79808b1b7921f3a765edb2b5bde54d53f75f2ff52ca72bc480af2f940e7ba923521e2a9f3d87cc3baaadbb1aff8be5b5ea1dd8cd13e0481fa2afd3d61e892082219f2b56302e0fca27f71b3915916eb598b1c6f89687c662bb4fc912d2f1c9527dec7f2985802e16b3fb45982
`define QX11 1032'h84d67a9d243ea4d7fa31629f471ba10a07c66598b80390f41c52cd01b01e9b93ca580bbb11ffc1769906adc9a56c28991128040b6476fda6adf11e8d329e02dfac964f171f79aa875a3518e9ccfd68aa73364dfc2d6751f38086c5e5539d0333bf6d4c003fca965dfd829db11edad2169d619ee4abb8e81e10c21b4dee7e5e075d
`define QY00 1032'h6aa7075afb6a9f8382d9f59f04868bde55d40d760da08b8f5dd685f44c79fd9650a1be993264612d690384068e3eb44ad7c2a52a3cc516af991b828aa8efcc8865b9b20111cd7faaa257920084d0e083b01e8871a3a0b2a402ce0e7438566b0d3773800e1568fd1a9961af7ee8c36fb8a16e41760461c6767541e1b891cd670177
`define QY01 1032'h656273d375b1dccf633ee6b4352d89cd2a35f50a9ba61865184b4593c156b6e4541a8046fda2da5d2bf194e5355898d54ac2339dc9cbc2e1ac8f711d8945edccb3ead62841ce77ad0e73bec1c81c0671dbd85cbffd7acf8634510a6e688714c92e9092297543c7a4b1d2cc2226dc4d13af5471d86d67710a13af95332c2d7c98ef
`define QY10 1032'h34b4f00004f6ec59d95112dfaa42a0fe500c3050972bed0de11d4ea99d009ab44ed5ee64818c1b093be37e509ab6f263451c41659355b9239cda55da46179b1671811c318ef1044473cf64bf80f1415eff58722564de026174e9a7af660cc25143d55e0ed4e0d2a42568ea096e5a3e8f715b359b33b3927a9df828250da37ab282
`define QY11 1032'h2e0d6129c895dd3b2a2e6fad425588723819e6e34620b57e67eed9e8532121415874438fdb1b10f99d39872cc37808bb38a93448e63ea57a7a5e6cb4715930c9ca36dc939ee61143269151e22a8f33ebf3901694ec00aee6f5f80411d5b9e43416314bed36f8ba3136c8d07b047147209aed63c1901caddee89e5813c50bfd3111
`define QY_00 1032'h5c0799f9933be2d12e3910bfadded44559f8cb7cfc020a2af23070becee7fbe01bd2921ca598fb82e0627e216564d01e1b8d12c774dbc61607fa4849a9241ddb14cb7bea4ea4762bee0b827e45e69bf38541d0e37ab3185b84b1f6f128a99752c86f2a7c953c585bbbf3a5cfc1e59047b3e73e89cb9e3989901374f218dd43a934
`define QY_01 1032'h614c2d8118f4a5854dd41faa7d37d6568596e3e86dfc7d5537bbb11f5a0b42921859d06eda5a82531d746d42be4aeb93a88d8453e7d519e3f48659b6c8cdfc96c69a57c31ea37e2981ef55bd029b76055987fc9520d8fb79532efaf6f878ed96d152186135618dd1a382892c83ccb2eca6010e2762988ef5f1a5c1777e7d2e11bc
`define QY_10 1032'h91f9b15489af95fad7c1f37f0822bf255fc0a8a27276a8ac6ee9a8097e615ec21d9e6251567141a70d8283d758ec9205ae33768c1e4b23a2043b74fa0bfc4f4d090411b9d180f1921c93afbf49c63b183607e72fb975c89e12965db5faf3400ebc0d4c7bd5c482d22fec6b453c4ec170e3fa4a649c4c6d85675d2e859d072ff829
`define QY_11 1032'h98a1402ac610a51986e496b1700fd7b177b2f20fc381e03be8181ccac840d83514000d25fce24bb6ac2c7afb302b7badbaa683a8cb62374b26b75e1fe0bab999b04e5157c18be49369d1c29ca028488b41d042c032531c18918801538b461e2be9b15e9d73ac9b451e8c84d3a637b8dfba681c3e3fe352211cb6fe96e59ead799a
`define TX00 1032'ha6956d27f52dc6f7460a7a97a5741f3b78d967e63f77a0b2e804e865e272cade37483ff1ccbf7092ded3f182434c3a528b123df309324a222d3df4d15f5fd0391d3f3a9b0458ebbabb62f0527fc93993d3cfa22c4ccb05e6a251512a9762a9b43ff301ba725bbb59639af50bd30865d6379700bbe99021736997d97deaa61a0288
`define TX01 1032'ha1e60a0f4df7a90eb30f2dc816893131194d296b2eb3c5479027ee25924d3dcb6ab2eb0bc380f1d7cf27c460b8eee6d62726c4b11344ba399fc7ff1ad487f5bbb7e632e2d44c019f69b8c692559c8cb28f4163c3119661f37b0cb22b13af8ada73cfc6fa132e20801dcb8ef907db5ed9a3f8b4312fb87070efb9461b84aa285bb2
`define TX10 1032'h1f842bd54a96d9a42b1d576b636d4ced5a61305ac79808b1b7921f3a765edb2b5bde54d53f75f2ff52ca72bc480af2f940e7ba923521e2a9f3d87cc3baaadbb1aff8be5b5ea1dd8cd13e0481fa2afd3d61e892082219f2b56302e0fca27f71b3915916eb598b1c6f89687c662bb4fc912d2f1c9527dec7f2985802e16b3fb45982
`define TX11 1032'h84d67a9d243ea4d7fa31629f471ba10a07c66598b80390f41c52cd01b01e9b93ca580bbb11ffc1769906adc9a56c28991128040b6476fda6adf11e8d329e02dfac964f171f79aa875a3518e9ccfd68aa73364dfc2d6751f38086c5e5539d0333bf6d4c003fca965dfd829db11edad2169d619ee4abb8e81e10c21b4dee7e5e075d
`define TY00 1032'h5c0799f9933be2d12e3910bfadded44559f8cb7cfc020a2af23070becee7fbe01bd2921ca598fb82e0627e216564d01e1b8d12c774dbc61607fa4849a9241ddb14cb7bea4ea4762bee0b827e45e69bf38541d0e37ab3185b84b1f6f128a99752c86f2a7c953c585bbbf3a5cfc1e59047b3e73e89cb9e3989901374f218dd43a934
`define TY01 1032'h614c2d8118f4a5854dd41faa7d37d6568596e3e86dfc7d5537bbb11f5a0b42921859d06eda5a82531d746d42be4aeb93a88d8453e7d519e3f48659b6c8cdfc96c69a57c31ea37e2981ef55bd029b76055987fc9520d8fb79532efaf6f878ed96d152186135618dd1a382892c83ccb2eca6010e2762988ef5f1a5c1777e7d2e11bc
`define TY10 1032'h91f9b15489af95fad7c1f37f0822bf255fc0a8a27276a8ac6ee9a8097e615ec21d9e6251567141a70d8283d758ec9205ae33768c1e4b23a2043b74fa0bfc4f4d090411b9d180f1921c93afbf49c63b183607e72fb975c89e12965db5faf3400ebc0d4c7bd5c482d22fec6b453c4ec170e3fa4a649c4c6d85675d2e859d072ff829
`define TY11 1032'h98a1402ac610a51986e496b1700fd7b177b2f20fc381e03be8181ccac840d83514000d25fce24bb6ac2c7afb302b7badbaa683a8cb62374b26b75e1fe0bab999b04e5157c18be49369d1c29ca028488b41d042c032531c18918801538b461e2be9b15e9d73ac9b451e8c84d3a637b8dfba681c3e3fe352211cb6fe96e59ead799a
`define TZ00 1032'h39515eab71597dab4eecf9a14d9a9fdc5033270cf65d6a45aff9094ce49e0689938baf4a2802a34fb699fdd80c5c7b970cb0480e4e5f233a5eea352badec159c857ad2149f8e0a296f9ceb8135488388ca9fa6aae1ac3500787ffa9a9efffda0001d5575555aaa89aaaaaab15556ffffaaaa80002ffffffffaaaa9555555555555
`define TZ01 1032'h0
`define TZ10 1032'h0
`define TZ11 1032'h0
