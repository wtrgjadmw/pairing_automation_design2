`define PX 461'hff7bd2bb2363911c351ef5d244fe7f56b026bfa6bca0b8539fb749787a6f2663784e39912ac1aa103307d1edb0325891e9f447494ff04cd4a73
`define PX_ 461'h55d9819a31721439703e736f04377c8041bc6de4f0298f5da8916ab213907f5e53b2b8d97e53addfd0f830125022fcc2c0b66376b01a5dd6038
`define PX3 461'h53c8cf86c07f68a954a20ef43c8f86562cade3dcdc4d99984e947414534e27a6d0e8c7de2e1a4e50911771c90fec5f0c6887805befbb9128a03
`define PY 461'h2f524ef3e7d4351e222708e3194309bb7e950f4361cc6aa157389e8e89709af50ba84b303e55327fd3061b98d6e92459594fe7a20aded355375
`define PY_ 461'h1260305616d0170378336605e2ff2f21b734e1e484afddd0ff110159c048f0accc058a73a6ac0257030f9e667296c30fb515ac31df52bd755736
`define QX0 461'h127721f8c7f8d061416ec7bf2436e4d9dc3ba9d0bc979f1ed2404bf9d610488ae5e0602e2cc9ef1ca4317eb837481ff2759c571b409e55ec8ab3`define QX1 461'h10988a5658d71b10402c3021e37bfbe656f77c1468e513d960a7ee0229991564ddbf57640c5b2435b5a3e1b27ae1fc6193b6ea482bca8a53c97a`define QY0 461'h469c6e4197a92e484947cfbcdabe6722732a97966873e5c5aedc3bc63b87151b76d5e9531b48d430e8a4557f09a6c3afb7b8ac11bea7f0eaaa5`define QY1 461'he63168650b4fba4ec163544f4d396aa20797c66450c5d02c22e7ce023b9c67096187453de96b0122c898dd8ea3e6c0da3d2e45df58e1160b05e`define QY_0 461'h10eb8e613bd2c770d5c1599846e7794b47eb895f5445661eb996c7864527890a6552b09178dcc83bf1b5bac80f6ae91a4f2f1feae4162b9c0006`define QY_1 461'h6f23ebf04985eb06e3fa14f1fbfc9134ea4b67275c0477852560e62852633eb86a79ad2cbfaa56cd3b6724715c6e947a6d7c64e0a729949fa4d`define TX0 461'h127721f8c7f8d061416ec7bf2436e4d9dc3ba9d0bc979f1ed2404bf9d610488ae5e0602e2cc9ef1ca4317eb837481ff2759c571b409e55ec8ab3`define TX1 461'h10988a5658d71b10402c3021e37bfbe656f77c1468e513d960a7ee0229991564ddbf57640c5b2435b5a3e1b27ae1fc6193b6ea482bca8a53c97a`define TY0 461'h10eb8e613bd2c770d5c1599846e7794b47eb895f5445661eb996c7864527890a6552b09178dcc83bf1b5bac80f6ae91a4f2f1feae4162b9c0006`define TY1 461'h6f23ebf04985eb06e3fa14f1fbfc9134ea4b67275c0477852560e62852633eb86a79ad2cbfaa56cd3b6724715c6e947a6d7c64e0a729949fa4d`define TZ0 461'haaaaabaaab2a5aaa5aa296beb6ca04290e1cd2745335b84eb7b74bd572005a3e33ff0d9556eaa80ffbfffdffffaaaaab5555553ffff55555555`define TZ1 461'h0