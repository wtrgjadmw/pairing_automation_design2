`define PX 440'h80389117112d1d884c9100144c38f7c7dd80c0d0da56b14030cb929b60f149188f5083df66b0db51c21ad22ba0bacd93993a236f5a0322
`define PX_ 440'h72c76eecbacb4c6407f7b65e991ae1b76150138db15aa1d0b0dc5ac23003a8855bc3276e62f72a7afc5390872ac01274661a873ca5a789
`define PX3 440'h8da9b341678eeeac912a49c9ff570dd859b16e140352c0afb0baca7491dee9abc2dde0506a6a8c2887e213d016b588b2cc59bfa20e5ebb
`define PY 440'h6aed5c7fbe224175bea7157bf4b288ebbb134019c96882e38a3bcef9e54d4169345b8c0590967bf731d964a37d84feac553bd917375d1f
`define PY_ 440'h8812a3840dd6287695e1a0f6f0a1509383bd9444c248d02d576c1e63aba7b034b6b81f48391189d58c94fe0f4df5e15baa18d194c84d8c
`define QX0 440'hbc935ba352b6ebc8c2289cd721e4322a2cd767950b1515d4a3550d2cd2ec1fa930b4a02671609df9c2ecb1458d41b97b86bc9388bcf261`define QX1 440'hddd42cd1ad6a742681cdb94f346243d4348956999d74f3fb23a9fd562e9183918f972db68d1fdbd4fb7b3270e5c86d8bc77ce9ea108eaf`define QY0 440'h5710e2faaf410247fb905205c1e49493342841dc4d4b45fb1355f276b913fa2332fb236b2476e75ddd54017f1913287300b1ffe33134ce`define QY1 440'hcc1285eecff53d8c24db4b96840479bed8c3a04de7044ee0da25ece9050092a98db8436e16c28535de46823c1bd81db9058333da489e16`define QY_0 440'h9bef1d091cb767a458f8646d236f44ec0aa892823e660d15ce51fae6d7e0f77ab81887e2a5311e6ee11a6133b267b794fea2aac8ce75dd`define QY_1 440'h26ed7a14fc032c602fad6adc614f5fc0660d3410a4ad0430078200748bf45ef45d5b67dfb2e58096e027e076afa2c24ef9d176d1b70c95`define TX0 440'hbc935ba352b6ebc8c2289cd721e4322a2cd767950b1515d4a3550d2cd2ec1fa930b4a02671609df9c2ecb1458d41b97b86bc9388bcf261`define TX1 440'hddd42cd1ad6a742681cdb94f346243d4348956999d74f3fb23a9fd562e9183918f972db68d1fdbd4fb7b3270e5c86d8bc77ce9ea108eaf`define TY0 440'h9bef1d091cb767a458f8646d236f44ec0aa892823e660d15ce51fae6d7e0f77ab81887e2a5311e6ee11a6133b267b794fea2aac8ce75dd`define TY1 440'h26ed7a14fc032c602fad6adc614f5fc0660d3410a4ad0430078200748bf45ef45d5b67dfb2e58096e027e076afa2c24ef9d176d1b70c95`define TZ0 440'hcfffffc34079613ab77498d1aac2680c12f2ba1744eacef1e5812a26f0b0e6214ec54b23657fa3341919d4d34851ff800ab5554005555`define TZ1 440'h0